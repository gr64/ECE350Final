module wallace_mult_32s(
	input[31:0] A, B,
	output[31:0] product, 
	//output[63:0] x, y,
	output overflow);
	
	wire a0_0, a0_1, a0_10, a0_11, a0_12, a0_13, a0_14, a0_15, a0_16, a0_17, a0_18, a0_19, a0_2, a0_20, a0_21, a0_22;
	wire a0_23, a0_24, a0_25, a0_26, a0_27, a0_28, a0_29, a0_3, a0_30, a0_31, a0_4, a0_5, a0_6, a0_7, a0_8, a0_9;
	wire a10_10, a10_11, a10_12, a10_13, a10_14, a10_15, a10_16, a10_17, a10_18, a10_19, a10_20, a10_21, a10_22, a10_23, a10_24, a10_25;
	wire a10_26, a10_27, a10_28, a10_29, a10_30, a10_31, a10_32, a10_33, a10_34, a10_35, a10_36, a10_37, a10_38, a10_39, a10_40, a10_41;
	wire a11_11, a11_12, a11_13, a11_14, a11_15, a11_16, a11_17, a11_18, a11_19, a11_20, a11_21, a11_22, a11_23, a11_24, a11_25, a11_26;
	wire a11_27, a11_28, a11_29, a11_30, a11_31, a11_32, a11_33, a11_34, a11_35, a11_36, a11_37, a11_38, a11_39, a11_40, a11_41, a11_42;
	wire a12_12, a12_13, a12_14, a12_15, a12_16, a12_17, a12_18, a12_19, a12_20, a12_21, a12_22, a12_23, a12_24, a12_25, a12_26, a12_27;
	wire a12_28, a12_29, a12_30, a12_31, a12_32, a12_33, a12_34, a12_35, a12_36, a12_37, a12_38, a12_39, a12_40, a12_41, a12_42, a12_43;
	wire a13_13, a13_14, a13_15, a13_16, a13_17, a13_18, a13_19, a13_20, a13_21, a13_22, a13_23, a13_24, a13_25, a13_26, a13_27, a13_28;
	wire a13_29, a13_30, a13_31, a13_32, a13_33, a13_34, a13_35, a13_36, a13_37, a13_38, a13_39, a13_40, a13_41, a13_42, a13_43, a13_44;
	wire a14_14, a14_15, a14_16, a14_17, a14_18, a14_19, a14_20, a14_21, a14_22, a14_23, a14_24, a14_25, a14_26, a14_27, a14_28, a14_29;
	wire a14_30, a14_31, a14_32, a14_33, a14_34, a14_35, a14_36, a14_37, a14_38, a14_39, a14_40, a14_41, a14_42, a14_43, a14_44, a14_45;
	wire a15_15, a15_16, a15_17, a15_18, a15_19, a15_20, a15_21, a15_22, a15_23, a15_24, a15_25, a15_26, a15_27, a15_28, a15_29, a15_30;
	wire a15_31, a15_32, a15_33, a15_34, a15_35, a15_36, a15_37, a15_38, a15_39, a15_40, a15_41, a15_42, a15_43, a15_44, a15_45, a15_46;
	wire a16_16, a16_17, a16_18, a16_19, a16_20, a16_21, a16_22, a16_23, a16_24, a16_25, a16_26, a16_27, a16_28, a16_29, a16_30, a16_31;
	wire a16_32, a16_33, a16_34, a16_35, a16_36, a16_37, a16_38, a16_39, a16_40, a16_41, a16_42, a16_43, a16_44, a16_45, a16_46, a16_47;
	wire a17_17, a17_18, a17_19, a17_20, a17_21, a17_22, a17_23, a17_24, a17_25, a17_26, a17_27, a17_28, a17_29, a17_30, a17_31, a17_32;
	wire a17_33, a17_34, a17_35, a17_36, a17_37, a17_38, a17_39, a17_40, a17_41, a17_42, a17_43, a17_44, a17_45, a17_46, a17_47, a17_48;
	wire a18_18, a18_19, a18_20, a18_21, a18_22, a18_23, a18_24, a18_25, a18_26, a18_27, a18_28, a18_29, a18_30, a18_31, a18_32, a18_33;
	wire a18_34, a18_35, a18_36, a18_37, a18_38, a18_39, a18_40, a18_41, a18_42, a18_43, a18_44, a18_45, a18_46, a18_47, a18_48, a18_49;
	wire a19_19, a19_20, a19_21, a19_22, a19_23, a19_24, a19_25, a19_26, a19_27, a19_28, a19_29, a19_30, a19_31, a19_32, a19_33, a19_34;
	wire a19_35, a19_36, a19_37, a19_38, a19_39, a19_40, a19_41, a19_42, a19_43, a19_44, a19_45, a19_46, a19_47, a19_48, a19_49, a19_50;
	wire a1_1, a1_10, a1_11, a1_12, a1_13, a1_14, a1_15, a1_16, a1_17, a1_18, a1_19, a1_2, a1_20, a1_21, a1_22, a1_23;
	wire a1_24, a1_25, a1_26, a1_27, a1_28, a1_29, a1_3, a1_30, a1_31, a1_32, a1_4, a1_5, a1_6, a1_7, a1_8, a1_9;
	wire a20_20, a20_21, a20_22, a20_23, a20_24, a20_25, a20_26, a20_27, a20_28, a20_29, a20_30, a20_31, a20_32, a20_33, a20_34, a20_35;
	wire a20_36, a20_37, a20_38, a20_39, a20_40, a20_41, a20_42, a20_43, a20_44, a20_45, a20_46, a20_47, a20_48, a20_49, a20_50, a20_51;
	wire a21_21, a21_22, a21_23, a21_24, a21_25, a21_26, a21_27, a21_28, a21_29, a21_30, a21_31, a21_32, a21_33, a21_34, a21_35, a21_36;
	wire a21_37, a21_38, a21_39, a21_40, a21_41, a21_42, a21_43, a21_44, a21_45, a21_46, a21_47, a21_48, a21_49, a21_50, a21_51, a21_52;
	wire a22_22, a22_23, a22_24, a22_25, a22_26, a22_27, a22_28, a22_29, a22_30, a22_31, a22_32, a22_33, a22_34, a22_35, a22_36, a22_37;
	wire a22_38, a22_39, a22_40, a22_41, a22_42, a22_43, a22_44, a22_45, a22_46, a22_47, a22_48, a22_49, a22_50, a22_51, a22_52, a22_53;
	wire a23_23, a23_24, a23_25, a23_26, a23_27, a23_28, a23_29, a23_30, a23_31, a23_32, a23_33, a23_34, a23_35, a23_36, a23_37, a23_38;
	wire a23_39, a23_40, a23_41, a23_42, a23_43, a23_44, a23_45, a23_46, a23_47, a23_48, a23_49, a23_50, a23_51, a23_52, a23_53, a23_54;
	wire a24_24, a24_25, a24_26, a24_27, a24_28, a24_29, a24_30, a24_31, a24_32, a24_33, a24_34, a24_35, a24_36, a24_37, a24_38, a24_39;
	wire a24_40, a24_41, a24_42, a24_43, a24_44, a24_45, a24_46, a24_47, a24_48, a24_49, a24_50, a24_51, a24_52, a24_53, a24_54, a24_55;
	wire a25_25, a25_26, a25_27, a25_28, a25_29, a25_30, a25_31, a25_32, a25_33, a25_34, a25_35, a25_36, a25_37, a25_38, a25_39, a25_40;
	wire a25_41, a25_42, a25_43, a25_44, a25_45, a25_46, a25_47, a25_48, a25_49, a25_50, a25_51, a25_52, a25_53, a25_54, a25_55, a25_56;
	wire a26_26, a26_27, a26_28, a26_29, a26_30, a26_31, a26_32, a26_33, a26_34, a26_35, a26_36, a26_37, a26_38, a26_39, a26_40, a26_41;
	wire a26_42, a26_43, a26_44, a26_45, a26_46, a26_47, a26_48, a26_49, a26_50, a26_51, a26_52, a26_53, a26_54, a26_55, a26_56, a26_57;
	wire a27_27, a27_28, a27_29, a27_30, a27_31, a27_32, a27_33, a27_34, a27_35, a27_36, a27_37, a27_38, a27_39, a27_40, a27_41, a27_42;
	wire a27_43, a27_44, a27_45, a27_46, a27_47, a27_48, a27_49, a27_50, a27_51, a27_52, a27_53, a27_54, a27_55, a27_56, a27_57, a27_58;
	wire a28_28, a28_29, a28_30, a28_31, a28_32, a28_33, a28_34, a28_35, a28_36, a28_37, a28_38, a28_39, a28_40, a28_41, a28_42, a28_43;
	wire a28_44, a28_45, a28_46, a28_47, a28_48, a28_49, a28_50, a28_51, a28_52, a28_53, a28_54, a28_55, a28_56, a28_57, a28_58, a28_59;
	wire a29_29, a29_30, a29_31, a29_32, a29_33, a29_34, a29_35, a29_36, a29_37, a29_38, a29_39, a29_40, a29_41, a29_42, a29_43, a29_44;
	wire a29_45, a29_46, a29_47, a29_48, a29_49, a29_50, a29_51, a29_52, a29_53, a29_54, a29_55, a29_56, a29_57, a29_58, a29_59, a29_60;
	wire a2_10, a2_11, a2_12, a2_13, a2_14, a2_15, a2_16, a2_17, a2_18, a2_19, a2_2, a2_20, a2_21, a2_22, a2_23, a2_24;
	wire a2_25, a2_26, a2_27, a2_28, a2_29, a2_3, a2_30, a2_31, a2_32, a2_33, a2_4, a2_5, a2_6, a2_7, a2_8, a2_9;
	wire a30_30, a30_31, a30_32, a30_33, a30_34, a30_35, a30_36, a30_37, a30_38, a30_39, a30_40, a30_41, a30_42, a30_43, a30_44, a30_45;
	wire a30_46, a30_47, a30_48, a30_49, a30_50, a30_51, a30_52, a30_53, a30_54, a30_55, a30_56, a30_57, a30_58, a30_59, a30_60, a30_61;
	wire a31_31, a31_32, a31_33, a31_34, a31_35, a31_36, a31_37, a31_38, a31_39, a31_40, a31_41, a31_42, a31_43, a31_44, a31_45, a31_46;
	wire a31_47, a31_48, a31_49, a31_50, a31_51, a31_52, a31_53, a31_54, a31_55, a31_56, a31_57, a31_58, a31_59, a31_60, a31_61, a31_62;
	wire a3_10, a3_11, a3_12, a3_13, a3_14, a3_15, a3_16, a3_17, a3_18, a3_19, a3_20, a3_21, a3_22, a3_23, a3_24, a3_25;
	wire a3_26, a3_27, a3_28, a3_29, a3_3, a3_30, a3_31, a3_32, a3_33, a3_34, a3_4, a3_5, a3_6, a3_7, a3_8, a3_9;
	wire a4_10, a4_11, a4_12, a4_13, a4_14, a4_15, a4_16, a4_17, a4_18, a4_19, a4_20, a4_21, a4_22, a4_23, a4_24, a4_25;
	wire a4_26, a4_27, a4_28, a4_29, a4_30, a4_31, a4_32, a4_33, a4_34, a4_35, a4_4, a4_5, a4_6, a4_7, a4_8, a4_9;
	wire a5_10, a5_11, a5_12, a5_13, a5_14, a5_15, a5_16, a5_17, a5_18, a5_19, a5_20, a5_21, a5_22, a5_23, a5_24, a5_25;
	wire a5_26, a5_27, a5_28, a5_29, a5_30, a5_31, a5_32, a5_33, a5_34, a5_35, a5_36, a5_5, a5_6, a5_7, a5_8, a5_9;
	wire a6_10, a6_11, a6_12, a6_13, a6_14, a6_15, a6_16, a6_17, a6_18, a6_19, a6_20, a6_21, a6_22, a6_23, a6_24, a6_25;
	wire a6_26, a6_27, a6_28, a6_29, a6_30, a6_31, a6_32, a6_33, a6_34, a6_35, a6_36, a6_37, a6_6, a6_7, a6_8, a6_9;
	wire a7_10, a7_11, a7_12, a7_13, a7_14, a7_15, a7_16, a7_17, a7_18, a7_19, a7_20, a7_21, a7_22, a7_23, a7_24, a7_25;
	wire a7_26, a7_27, a7_28, a7_29, a7_30, a7_31, a7_32, a7_33, a7_34, a7_35, a7_36, a7_37, a7_38, a7_7, a7_8, a7_9;
	wire a8_10, a8_11, a8_12, a8_13, a8_14, a8_15, a8_16, a8_17, a8_18, a8_19, a8_20, a8_21, a8_22, a8_23, a8_24, a8_25;
	wire a8_26, a8_27, a8_28, a8_29, a8_30, a8_31, a8_32, a8_33, a8_34, a8_35, a8_36, a8_37, a8_38, a8_39, a8_8, a8_9;
	wire a9_10, a9_11, a9_12, a9_13, a9_14, a9_15, a9_16, a9_17, a9_18, a9_19, a9_20, a9_21, a9_22, a9_23, a9_24, a9_25;
	wire a9_26, a9_27, a9_28, a9_29, a9_30, a9_31, a9_32, a9_33, a9_34, a9_35, a9_36, a9_37, a9_38, a9_39, a9_40, a9_9;
	wire ap0_31, ap10_41, ap11_42, ap12_43, ap13_44, ap14_45, ap15_46, ap16_47, ap17_48, ap18_49, ap19_50, ap1_32, ap20_51, ap21_52, ap22_53, ap23_54;
	wire ap24_55, ap25_56, ap26_57, ap27_58, ap28_59, ap29_60, ap2_33, ap30_61, ap31_31, ap31_32, ap31_33, ap31_34, ap31_35, ap31_36, ap31_37, ap31_38;
	wire ap31_39, ap31_40, ap31_41, ap31_42, ap31_43, ap31_44, ap31_45, ap31_46, ap31_47, ap31_48, ap31_49, ap31_50, ap31_51, ap31_52, ap31_53, ap31_54;
	wire ap31_55, ap31_56, ap31_57, ap31_58, ap31_59, ap31_60, ap31_61, ap3_34, ap4_35, ap5_36, ap6_37, ap7_38, ap8_39, ap9_40, c10_0_0, c10_0_1;
	wire c10_0_2, c10_0_3, c10_1_0, c10_1_1, c10_2_0, c10_2_1, c10_3_0, c10_4_0, c10_5_0, c10_6_0, c10_7_0, c11_0_0, c11_0_1, c11_0_2, c11_0_3, c11_1_0;
	wire c11_1_1, c11_1_2, c11_2_0, c11_2_1, c11_3_0, c11_4_0, c11_5_0, c11_6_0, c11_7_0, c12_0_0, c12_0_1, c12_0_2, c12_0_3, c12_1_0, c12_1_1, c12_1_2;
	wire c12_2_0, c12_2_1, c12_3_0, c12_4_0, c12_5_0, c12_6_0, c12_7_0, c13_0_0, c13_0_1, c13_0_2, c13_0_3, c13_0_4, c13_1_0, c13_1_1, c13_1_2, c13_2_0;
	wire c13_2_1, c13_3_0, c13_4_0, c13_5_0, c13_6_0, c13_7_0, c14_0_0, c14_0_1, c14_0_2, c14_0_3, c14_0_4, c14_1_0, c14_1_1, c14_1_2, c14_2_0, c14_2_1;
	wire c14_3_0, c14_3_1, c14_4_0, c14_5_0, c14_6_0, c14_7_0, c15_0_0, c15_0_1, c15_0_2, c15_0_3, c15_0_4, c15_1_0, c15_1_1, c15_1_2, c15_1_3, c15_2_0;
	wire c15_2_1, c15_3_0, c15_3_1, c15_4_0, c15_5_0, c15_6_0, c15_7_0, c16_0_0, c16_0_1, c16_0_2, c16_0_3, c16_0_4, c16_0_5, c16_1_0, c16_1_1, c16_1_2;
	wire c16_1_3, c16_2_0, c16_2_1, c16_2_2, c16_3_0, c16_3_1, c16_4_0, c16_5_0, c16_6_0, c16_7_0, c17_0_0, c17_0_1, c17_0_2, c17_0_3, c17_0_4, c17_0_5;
	wire c17_1_0, c17_1_1, c17_1_2, c17_1_3, c17_2_0, c17_2_1, c17_2_2, c17_3_0, c17_3_1, c17_4_0, c17_5_0, c17_6_0, c17_7_0, c18_0_0, c18_0_1, c18_0_2;
	wire c18_0_3, c18_0_4, c18_0_5, c18_1_0, c18_1_1, c18_1_2, c18_1_3, c18_2_0, c18_2_1, c18_2_2, c18_3_0, c18_3_1, c18_4_0, c18_5_0, c18_6_0, c18_7_0;
	wire c19_0_0, c19_0_1, c19_0_2, c19_0_3, c19_0_4, c19_0_5, c19_0_6, c19_1_0, c19_1_1, c19_1_2, c19_1_3, c19_2_0, c19_2_1, c19_2_2, c19_3_0, c19_3_1;
	wire c19_4_0, c19_5_0, c19_6_0, c19_7_0, c1_0_0, c20_0_0, c20_0_1, c20_0_2, c20_0_3, c20_0_4, c20_0_5, c20_0_6, c20_1_0, c20_1_1, c20_1_2, c20_1_3;
	wire c20_1_4, c20_2_0, c20_2_1, c20_2_2, c20_3_0, c20_3_1, c20_4_0, c20_5_0, c20_6_0, c20_7_0, c21_0_0, c21_0_1, c21_0_2, c21_0_3, c21_0_4, c21_0_5;
	wire c21_0_6, c21_1_0, c21_1_1, c21_1_2, c21_1_3, c21_1_4, c21_2_0, c21_2_1, c21_2_2, c21_3_0, c21_3_1, c21_4_0, c21_4_1, c21_5_0, c21_6_0, c21_7_0;
	wire c22_0_0, c22_0_1, c22_0_2, c22_0_3, c22_0_4, c22_0_5, c22_0_6, c22_0_7, c22_1_0, c22_1_1, c22_1_2, c22_1_3, c22_1_4, c22_2_0, c22_2_1, c22_2_2;
	wire c22_3_0, c22_3_1, c22_4_0, c22_4_1, c22_5_0, c22_6_0, c22_7_0, c23_0_0, c23_0_1, c23_0_2, c23_0_3, c23_0_4, c23_0_5, c23_0_6, c23_0_7, c23_1_0;
	wire c23_1_1, c23_1_2, c23_1_3, c23_1_4, c23_2_0, c23_2_1, c23_2_2, c23_2_3, c23_3_0, c23_3_1, c23_4_0, c23_4_1, c23_5_0, c23_6_0, c23_7_0, c24_0_0;
	wire c24_0_1, c24_0_2, c24_0_3, c24_0_4, c24_0_5, c24_0_6, c24_0_7, c24_1_0, c24_1_1, c24_1_2, c24_1_3, c24_1_4, c24_1_5, c24_2_0, c24_2_1, c24_2_2;
	wire c24_2_3, c24_3_0, c24_3_1, c24_3_2, c24_4_0, c24_4_1, c24_5_0, c24_6_0, c24_7_0, c25_0_0, c25_0_1, c25_0_2, c25_0_3, c25_0_4, c25_0_5, c25_0_6;
	wire c25_0_7, c25_0_8, c25_1_0, c25_1_1, c25_1_2, c25_1_3, c25_1_4, c25_1_5, c25_2_0, c25_2_1, c25_2_2, c25_2_3, c25_3_0, c25_3_1, c25_3_2, c25_4_0;
	wire c25_4_1, c25_5_0, c25_6_0, c25_7_0, c26_0_0, c26_0_1, c26_0_2, c26_0_3, c26_0_4, c26_0_5, c26_0_6, c26_0_7, c26_0_8, c26_1_0, c26_1_1, c26_1_2;
	wire c26_1_3, c26_1_4, c26_1_5, c26_2_0, c26_2_1, c26_2_2, c26_2_3, c26_3_0, c26_3_1, c26_3_2, c26_4_0, c26_4_1, c26_5_0, c26_6_0, c26_7_0, c27_0_0;
	wire c27_0_1, c27_0_2, c27_0_3, c27_0_4, c27_0_5, c27_0_6, c27_0_7, c27_0_8, c27_1_0, c27_1_1, c27_1_2, c27_1_3, c27_1_4, c27_1_5, c27_2_0, c27_2_1;
	wire c27_2_2, c27_2_3, c27_3_0, c27_3_1, c27_3_2, c27_4_0, c27_4_1, c27_5_0, c27_6_0, c27_7_0, c28_0_0, c28_0_1, c28_0_2, c28_0_3, c28_0_4, c28_0_5;
	wire c28_0_6, c28_0_7, c28_0_8, c28_0_9, c28_1_0, c28_1_1, c28_1_2, c28_1_3, c28_1_4, c28_1_5, c28_2_0, c28_2_1, c28_2_2, c28_2_3, c28_3_0, c28_3_1;
	wire c28_3_2, c28_4_0, c28_4_1, c28_5_0, c28_6_0, c28_7_0, c29_0_0, c29_0_1, c29_0_2, c29_0_3, c29_0_4, c29_0_5, c29_0_6, c29_0_7, c29_0_8, c29_0_9;
	wire c29_1_0, c29_1_1, c29_1_2, c29_1_3, c29_1_4, c29_1_5, c29_1_6, c29_2_0, c29_2_1, c29_2_2, c29_2_3, c29_3_0, c29_3_1, c29_3_2, c29_4_0, c29_4_1;
	wire c29_5_0, c29_6_0, c29_7_0, c2_0_0, c2_1_0, c30_0_0, c30_0_1, c30_0_2, c30_0_3, c30_0_4, c30_0_5, c30_0_6, c30_0_7, c30_0_8, c30_0_9, c30_1_0;
	wire c30_1_1, c30_1_2, c30_1_3, c30_1_4, c30_1_5, c30_1_6, c30_2_0, c30_2_1, c30_2_2, c30_2_3, c30_2_4, c30_3_0, c30_3_1, c30_3_2, c30_4_0, c30_4_1;
	wire c30_5_0, c30_6_0, c30_7_0, c31_0_0, c31_0_1, c31_0_10, c31_0_2, c31_0_3, c31_0_4, c31_0_5, c31_0_6, c31_0_7, c31_0_8, c31_0_9, c31_1_0, c31_1_1;
	wire c31_1_2, c31_1_3, c31_1_4, c31_1_5, c31_1_6, c31_2_0, c31_2_1, c31_2_2, c31_2_3, c31_2_4, c31_3_0, c31_3_1, c31_3_2, c31_4_0, c31_4_1, c31_5_0;
	wire c31_5_1, c31_6_0, c31_7_0, c32_0_0, c32_0_1, c32_0_10, c32_0_2, c32_0_3, c32_0_4, c32_0_5, c32_0_6, c32_0_7, c32_0_8, c32_0_9, c32_1_0, c32_1_1;
	wire c32_1_2, c32_1_3, c32_1_4, c32_1_5, c32_1_6, c32_2_0, c32_2_1, c32_2_2, c32_2_3, c32_2_4, c32_3_0, c32_3_1, c32_3_2, c32_4_0, c32_4_1, c32_5_0;
	wire c32_5_1, c32_6_0, c32_7_0, c33_0_0, c33_0_1, c33_0_2, c33_0_3, c33_0_4, c33_0_5, c33_0_6, c33_0_7, c33_0_8, c33_0_9, c33_1_0, c33_1_1, c33_1_2;
	wire c33_1_3, c33_1_4, c33_1_5, c33_1_6, c33_2_0, c33_2_1, c33_2_2, c33_2_3, c33_2_4, c33_3_0, c33_3_1, c33_3_2, c33_4_0, c33_4_1, c33_5_0, c33_5_1;
	wire c33_6_0, c33_7_0, c34_0_0, c34_0_1, c34_0_2, c34_0_3, c34_0_4, c34_0_5, c34_0_6, c34_0_7, c34_0_8, c34_0_9, c34_1_0, c34_1_1, c34_1_2, c34_1_3;
	wire c34_1_4, c34_1_5, c34_1_6, c34_2_0, c34_2_1, c34_2_2, c34_2_3, c34_2_4, c34_3_0, c34_3_1, c34_3_2, c34_4_0, c34_4_1, c34_5_0, c34_5_1, c34_6_0;
	wire c34_7_0, c35_0_0, c35_0_1, c35_0_2, c35_0_3, c35_0_4, c35_0_5, c35_0_6, c35_0_7, c35_0_8, c35_1_0, c35_1_1, c35_1_2, c35_1_3, c35_1_4, c35_1_5;
	wire c35_1_6, c35_2_0, c35_2_1, c35_2_2, c35_2_3, c35_2_4, c35_3_0, c35_3_1, c35_3_2, c35_4_0, c35_4_1, c35_5_0, c35_5_1, c35_6_0, c35_7_0, c36_0_0;
	wire c36_0_1, c36_0_2, c36_0_3, c36_0_4, c36_0_5, c36_0_6, c36_0_7, c36_0_8, c36_1_0, c36_1_1, c36_1_2, c36_1_3, c36_1_4, c36_1_5, c36_2_0, c36_2_1;
	wire c36_2_2, c36_2_3, c36_3_0, c36_3_1, c36_3_2, c36_4_0, c36_4_1, c36_5_0, c36_5_1, c36_6_0, c36_7_0, c37_0_0, c37_0_1, c37_0_2, c37_0_3, c37_0_4;
	wire c37_0_5, c37_0_6, c37_0_7, c37_0_8, c37_1_0, c37_1_1, c37_1_2, c37_1_3, c37_1_4, c37_1_5, c37_2_0, c37_2_1, c37_2_2, c37_2_3, c37_3_0, c37_3_1;
	wire c37_3_2, c37_4_0, c37_4_1, c37_5_0, c37_6_0, c37_7_0, c38_0_0, c38_0_1, c38_0_2, c38_0_3, c38_0_4, c38_0_5, c38_0_6, c38_0_7, c38_1_0, c38_1_1;
	wire c38_1_2, c38_1_3, c38_1_4, c38_1_5, c38_2_0, c38_2_1, c38_2_2, c38_2_3, c38_3_0, c38_3_1, c38_3_2, c38_4_0, c38_4_1, c38_5_0, c38_6_0, c38_7_0;
	wire c39_0_0, c39_0_1, c39_0_2, c39_0_3, c39_0_4, c39_0_5, c39_0_6, c39_0_7, c39_1_0, c39_1_1, c39_1_2, c39_1_3, c39_1_4, c39_2_0, c39_2_1, c39_2_2;
	wire c39_2_3, c39_3_0, c39_3_1, c39_3_2, c39_4_0, c39_4_1, c39_5_0, c39_6_0, c39_7_0, c3_0_0, c3_1_0, c3_2_0, c40_0_0, c40_0_1, c40_0_2, c40_0_3;
	wire c40_0_4, c40_0_5, c40_0_6, c40_0_7, c40_1_0, c40_1_1, c40_1_2, c40_1_3, c40_1_4, c40_2_0, c40_2_1, c40_2_2, c40_2_3, c40_3_0, c40_3_1, c40_3_2;
	wire c40_4_0, c40_4_1, c40_5_0, c40_6_0, c40_7_0, c41_0_0, c41_0_1, c41_0_2, c41_0_3, c41_0_4, c41_0_5, c41_0_6, c41_1_0, c41_1_1, c41_1_2, c41_1_3;
	wire c41_1_4, c41_2_0, c41_2_1, c41_2_2, c41_2_3, c41_3_0, c41_3_1, c41_3_2, c41_4_0, c41_4_1, c41_5_0, c41_6_0, c41_7_0, c42_0_0, c42_0_1, c42_0_2;
	wire c42_0_3, c42_0_4, c42_0_5, c42_0_6, c42_1_0, c42_1_1, c42_1_2, c42_1_3, c42_1_4, c42_2_0, c42_2_1, c42_2_2, c42_3_0, c42_3_1, c42_3_2, c42_4_0;
	wire c42_4_1, c42_5_0, c42_6_0, c42_7_0, c43_0_0, c43_0_1, c43_0_2, c43_0_3, c43_0_4, c43_0_5, c43_0_6, c43_1_0, c43_1_1, c43_1_2, c43_1_3, c43_1_4;
	wire c43_2_0, c43_2_1, c43_2_2, c43_3_0, c43_3_1, c43_4_0, c43_4_1, c43_5_0, c43_6_0, c43_7_0, c44_0_0, c44_0_1, c44_0_2, c44_0_3, c44_0_4, c44_0_5;
	wire c44_1_0, c44_1_1, c44_1_2, c44_1_3, c44_1_4, c44_2_0, c44_2_1, c44_2_2, c44_3_0, c44_3_1, c44_4_0, c44_4_1, c44_5_0, c44_6_0, c44_7_0, c45_0_0;
	wire c45_0_1, c45_0_2, c45_0_3, c45_0_4, c45_0_5, c45_1_0, c45_1_1, c45_1_2, c45_1_3, c45_2_0, c45_2_1, c45_2_2, c45_3_0, c45_3_1, c45_4_0, c45_5_0;
	wire c45_6_0, c45_7_0, c46_0_0, c46_0_1, c46_0_2, c46_0_3, c46_0_4, c46_0_5, c46_1_0, c46_1_1, c46_1_2, c46_1_3, c46_2_0, c46_2_1, c46_2_2, c46_3_0;
	wire c46_3_1, c46_4_0, c46_5_0, c46_6_0, c46_7_0, c47_0_0, c47_0_1, c47_0_2, c47_0_3, c47_0_4, c47_1_0, c47_1_1, c47_1_2, c47_1_3, c47_2_0, c47_2_1;
	wire c47_2_2, c47_3_0, c47_3_1, c47_4_0, c47_5_0, c47_6_0, c47_7_0, c48_0_0, c48_0_1, c48_0_2, c48_0_3, c48_0_4, c48_1_0, c48_1_1, c48_1_2, c48_2_0;
	wire c48_2_1, c48_2_2, c48_3_0, c48_3_1, c48_4_0, c48_5_0, c48_6_0, c48_7_0, c49_0_0, c49_0_1, c49_0_2, c49_0_3, c49_0_4, c49_1_0, c49_1_1, c49_1_2;
	wire c49_2_0, c49_2_1, c49_3_0, c49_3_1, c49_4_0, c49_5_0, c49_6_0, c49_7_0, c4_0_0, c4_0_1, c4_1_0, c4_2_0, c4_3_0, c50_0_0, c50_0_1, c50_0_2;
	wire c50_0_3, c50_1_0, c50_1_1, c50_1_2, c50_2_0, c50_2_1, c50_3_0, c50_3_1, c50_4_0, c50_5_0, c50_6_0, c50_7_0, c51_0_0, c51_0_1, c51_0_2, c51_0_3;
	wire c51_1_0, c51_1_1, c51_1_2, c51_2_0, c51_2_1, c51_3_0, c51_4_0, c51_5_0, c51_6_0, c51_7_0, c52_0_0, c52_0_1, c52_0_2, c52_0_3, c52_1_0, c52_1_1;
	wire c52_1_2, c52_2_0, c52_2_1, c52_3_0, c52_4_0, c52_5_0, c52_6_0, c52_7_0, c53_0_0, c53_0_1, c53_0_2, c53_1_0, c53_1_1, c53_1_2, c53_2_0, c53_2_1;
	wire c53_3_0, c53_4_0, c53_5_0, c53_6_0, c53_7_0, c54_0_0, c54_0_1, c54_0_2, c54_1_0, c54_1_1, c54_2_0, c54_2_1, c54_3_0, c54_4_0, c54_5_0, c54_6_0;
	wire c54_7_0, c55_0_0, c55_0_1, c55_0_2, c55_1_0, c55_1_1, c55_2_0, c55_3_0, c55_4_0, c55_5_0, c55_6_0, c55_7_0, c56_0_0, c56_0_1, c56_1_0, c56_1_1;
	wire c56_2_0, c56_3_0, c56_4_0, c56_5_0, c56_6_0, c56_7_0, c57_0_0, c57_0_1, c57_1_0, c57_2_0, c57_3_0, c57_4_0, c57_5_0, c57_6_0, c57_7_0, c58_0_0;
	wire c58_0_1, c58_1_0, c58_2_0, c58_3_0, c58_4_0, c58_5_0, c58_6_0, c58_7_0, c59_0_0, c59_1_0, c59_2_0, c59_3_0, c59_4_0, c59_5_0, c59_6_0, c59_7_0;
	wire c5_0_0, c5_0_1, c5_1_0, c5_2_0, c5_3_0, c5_4_0, c60_0_0, c60_1_0, c60_2_0, c60_3_0, c60_4_0, c60_5_0, c60_6_0, c60_7_0, c61_0_0, c61_1_0;
	wire c61_2_0, c61_3_0, c61_4_0, c61_5_0, c61_6_0, c61_7_0, c62_1_0, c62_2_0, c62_3_0, c62_4_0, c62_5_0, c62_6_0, c62_7_0, c63_2_0, c63_3_0, c63_4_0;
	wire c63_5_0, c63_6_0, c63_7_0, c6_0_0, c6_0_1, c6_1_0, c6_1_1, c6_2_0, c6_3_0, c6_4_0, c6_5_0, c7_0_0, c7_0_1, c7_0_2, c7_1_0, c7_1_1;
	wire c7_2_0, c7_3_0, c7_4_0, c7_5_0, c7_6_0, c8_0_0, c8_0_1, c8_0_2, c8_1_0, c8_1_1, c8_2_0, c8_3_0, c8_4_0, c8_5_0, c8_6_0, c8_7_0;
	wire c9_0_0, c9_0_1, c9_0_2, c9_1_0, c9_1_1, c9_2_0, c9_2_1, c9_3_0, c9_4_0, c9_5_0, c9_6_0, c9_7_0, s10_0_0, s10_0_1, s10_0_2, s10_0_3;
	wire s10_1_0, s10_1_1, s10_2_0, s10_2_1, s10_3_0, s10_4_0, s10_5_0, s10_6_0, s10_7_0, s11_0_0, s11_0_1, s11_0_2, s11_0_3, s11_1_0, s11_1_1, s11_1_2;
	wire s11_2_0, s11_2_1, s11_3_0, s11_4_0, s11_5_0, s11_6_0, s11_7_0, s12_0_0, s12_0_1, s12_0_2, s12_0_3, s12_1_0, s12_1_1, s12_1_2, s12_2_0, s12_2_1;
	wire s12_3_0, s12_4_0, s12_5_0, s12_6_0, s12_7_0, s13_0_0, s13_0_1, s13_0_2, s13_0_3, s13_0_4, s13_1_0, s13_1_1, s13_1_2, s13_2_0, s13_2_1, s13_3_0;
	wire s13_4_0, s13_5_0, s13_6_0, s13_7_0, s14_0_0, s14_0_1, s14_0_2, s14_0_3, s14_0_4, s14_1_0, s14_1_1, s14_1_2, s14_2_0, s14_2_1, s14_3_0, s14_3_1;
	wire s14_4_0, s14_5_0, s14_6_0, s14_7_0, s15_0_0, s15_0_1, s15_0_2, s15_0_3, s15_0_4, s15_1_0, s15_1_1, s15_1_2, s15_1_3, s15_2_0, s15_2_1, s15_3_0;
	wire s15_3_1, s15_4_0, s15_5_0, s15_6_0, s15_7_0, s16_0_0, s16_0_1, s16_0_2, s16_0_3, s16_0_4, s16_0_5, s16_1_0, s16_1_1, s16_1_2, s16_1_3, s16_2_0;
	wire s16_2_1, s16_2_2, s16_3_0, s16_3_1, s16_4_0, s16_5_0, s16_6_0, s16_7_0, s17_0_0, s17_0_1, s17_0_2, s17_0_3, s17_0_4, s17_0_5, s17_1_0, s17_1_1;
	wire s17_1_2, s17_1_3, s17_2_0, s17_2_1, s17_2_2, s17_3_0, s17_3_1, s17_4_0, s17_5_0, s17_6_0, s17_7_0, s18_0_0, s18_0_1, s18_0_2, s18_0_3, s18_0_4;
	wire s18_0_5, s18_1_0, s18_1_1, s18_1_2, s18_1_3, s18_2_0, s18_2_1, s18_2_2, s18_3_0, s18_3_1, s18_4_0, s18_5_0, s18_6_0, s18_7_0, s19_0_0, s19_0_1;
	wire s19_0_2, s19_0_3, s19_0_4, s19_0_5, s19_0_6, s19_1_0, s19_1_1, s19_1_2, s19_1_3, s19_2_0, s19_2_1, s19_2_2, s19_3_0, s19_3_1, s19_4_0, s19_5_0;
	wire s19_6_0, s19_7_0, s1_0_0, s20_0_0, s20_0_1, s20_0_2, s20_0_3, s20_0_4, s20_0_5, s20_0_6, s20_1_0, s20_1_1, s20_1_2, s20_1_3, s20_1_4, s20_2_0;
	wire s20_2_1, s20_2_2, s20_3_0, s20_3_1, s20_4_0, s20_5_0, s20_6_0, s20_7_0, s21_0_0, s21_0_1, s21_0_2, s21_0_3, s21_0_4, s21_0_5, s21_0_6, s21_1_0;
	wire s21_1_1, s21_1_2, s21_1_3, s21_1_4, s21_2_0, s21_2_1, s21_2_2, s21_3_0, s21_3_1, s21_4_0, s21_4_1, s21_5_0, s21_6_0, s21_7_0, s22_0_0, s22_0_1;
	wire s22_0_2, s22_0_3, s22_0_4, s22_0_5, s22_0_6, s22_0_7, s22_1_0, s22_1_1, s22_1_2, s22_1_3, s22_1_4, s22_2_0, s22_2_1, s22_2_2, s22_3_0, s22_3_1;
	wire s22_4_0, s22_4_1, s22_5_0, s22_6_0, s22_7_0, s23_0_0, s23_0_1, s23_0_2, s23_0_3, s23_0_4, s23_0_5, s23_0_6, s23_0_7, s23_1_0, s23_1_1, s23_1_2;
	wire s23_1_3, s23_1_4, s23_2_0, s23_2_1, s23_2_2, s23_2_3, s23_3_0, s23_3_1, s23_4_0, s23_4_1, s23_5_0, s23_6_0, s23_7_0, s24_0_0, s24_0_1, s24_0_2;
	wire s24_0_3, s24_0_4, s24_0_5, s24_0_6, s24_0_7, s24_1_0, s24_1_1, s24_1_2, s24_1_3, s24_1_4, s24_1_5, s24_2_0, s24_2_1, s24_2_2, s24_2_3, s24_3_0;
	wire s24_3_1, s24_3_2, s24_4_0, s24_4_1, s24_5_0, s24_6_0, s24_7_0, s25_0_0, s25_0_1, s25_0_2, s25_0_3, s25_0_4, s25_0_5, s25_0_6, s25_0_7, s25_0_8;
	wire s25_1_0, s25_1_1, s25_1_2, s25_1_3, s25_1_4, s25_1_5, s25_2_0, s25_2_1, s25_2_2, s25_2_3, s25_3_0, s25_3_1, s25_3_2, s25_4_0, s25_4_1, s25_5_0;
	wire s25_6_0, s25_7_0, s26_0_0, s26_0_1, s26_0_2, s26_0_3, s26_0_4, s26_0_5, s26_0_6, s26_0_7, s26_0_8, s26_1_0, s26_1_1, s26_1_2, s26_1_3, s26_1_4;
	wire s26_1_5, s26_2_0, s26_2_1, s26_2_2, s26_2_3, s26_3_0, s26_3_1, s26_3_2, s26_4_0, s26_4_1, s26_5_0, s26_6_0, s26_7_0, s27_0_0, s27_0_1, s27_0_2;
	wire s27_0_3, s27_0_4, s27_0_5, s27_0_6, s27_0_7, s27_0_8, s27_1_0, s27_1_1, s27_1_2, s27_1_3, s27_1_4, s27_1_5, s27_2_0, s27_2_1, s27_2_2, s27_2_3;
	wire s27_3_0, s27_3_1, s27_3_2, s27_4_0, s27_4_1, s27_5_0, s27_6_0, s27_7_0, s28_0_0, s28_0_1, s28_0_2, s28_0_3, s28_0_4, s28_0_5, s28_0_6, s28_0_7;
	wire s28_0_8, s28_0_9, s28_1_0, s28_1_1, s28_1_2, s28_1_3, s28_1_4, s28_1_5, s28_2_0, s28_2_1, s28_2_2, s28_2_3, s28_3_0, s28_3_1, s28_3_2, s28_4_0;
	wire s28_4_1, s28_5_0, s28_6_0, s28_7_0, s29_0_0, s29_0_1, s29_0_2, s29_0_3, s29_0_4, s29_0_5, s29_0_6, s29_0_7, s29_0_8, s29_0_9, s29_1_0, s29_1_1;
	wire s29_1_2, s29_1_3, s29_1_4, s29_1_5, s29_1_6, s29_2_0, s29_2_1, s29_2_2, s29_2_3, s29_3_0, s29_3_1, s29_3_2, s29_4_0, s29_4_1, s29_5_0, s29_6_0;
	wire s29_7_0, s2_0_0, s2_1_0, s30_0_0, s30_0_1, s30_0_2, s30_0_3, s30_0_4, s30_0_5, s30_0_6, s30_0_7, s30_0_8, s30_0_9, s30_1_0, s30_1_1, s30_1_2;
	wire s30_1_3, s30_1_4, s30_1_5, s30_1_6, s30_2_0, s30_2_1, s30_2_2, s30_2_3, s30_2_4, s30_3_0, s30_3_1, s30_3_2, s30_4_0, s30_4_1, s30_5_0, s30_6_0;
	wire s30_7_0, s31_0_0, s31_0_1, s31_0_10, s31_0_2, s31_0_3, s31_0_4, s31_0_5, s31_0_6, s31_0_7, s31_0_8, s31_0_9, s31_1_0, s31_1_1, s31_1_2, s31_1_3;
	wire s31_1_4, s31_1_5, s31_1_6, s31_2_0, s31_2_1, s31_2_2, s31_2_3, s31_2_4, s31_3_0, s31_3_1, s31_3_2, s31_4_0, s31_4_1, s31_5_0, s31_5_1, s31_6_0;
	wire s31_7_0, s32_0_0, s32_0_1, s32_0_10, s32_0_2, s32_0_3, s32_0_4, s32_0_5, s32_0_6, s32_0_7, s32_0_8, s32_0_9, s32_1_0, s32_1_1, s32_1_2, s32_1_3;
	wire s32_1_4, s32_1_5, s32_1_6, s32_2_0, s32_2_1, s32_2_2, s32_2_3, s32_2_4, s32_3_0, s32_3_1, s32_3_2, s32_4_0, s32_4_1, s32_5_0, s32_5_1, s32_6_0;
	wire s32_7_0, s33_0_0, s33_0_1, s33_0_2, s33_0_3, s33_0_4, s33_0_5, s33_0_6, s33_0_7, s33_0_8, s33_0_9, s33_1_0, s33_1_1, s33_1_2, s33_1_3, s33_1_4;
	wire s33_1_5, s33_1_6, s33_2_0, s33_2_1, s33_2_2, s33_2_3, s33_2_4, s33_3_0, s33_3_1, s33_3_2, s33_4_0, s33_4_1, s33_5_0, s33_5_1, s33_6_0, s33_7_0;
	wire s34_0_0, s34_0_1, s34_0_2, s34_0_3, s34_0_4, s34_0_5, s34_0_6, s34_0_7, s34_0_8, s34_0_9, s34_1_0, s34_1_1, s34_1_2, s34_1_3, s34_1_4, s34_1_5;
	wire s34_1_6, s34_2_0, s34_2_1, s34_2_2, s34_2_3, s34_2_4, s34_3_0, s34_3_1, s34_3_2, s34_4_0, s34_4_1, s34_5_0, s34_5_1, s34_6_0, s34_7_0, s35_0_0;
	wire s35_0_1, s35_0_2, s35_0_3, s35_0_4, s35_0_5, s35_0_6, s35_0_7, s35_0_8, s35_1_0, s35_1_1, s35_1_2, s35_1_3, s35_1_4, s35_1_5, s35_1_6, s35_2_0;
	wire s35_2_1, s35_2_2, s35_2_3, s35_2_4, s35_3_0, s35_3_1, s35_3_2, s35_4_0, s35_4_1, s35_5_0, s35_5_1, s35_6_0, s35_7_0, s36_0_0, s36_0_1, s36_0_2;
	wire s36_0_3, s36_0_4, s36_0_5, s36_0_6, s36_0_7, s36_0_8, s36_1_0, s36_1_1, s36_1_2, s36_1_3, s36_1_4, s36_1_5, s36_2_0, s36_2_1, s36_2_2, s36_2_3;
	wire s36_3_0, s36_3_1, s36_3_2, s36_4_0, s36_4_1, s36_5_0, s36_5_1, s36_6_0, s36_7_0, s37_0_0, s37_0_1, s37_0_2, s37_0_3, s37_0_4, s37_0_5, s37_0_6;
	wire s37_0_7, s37_0_8, s37_1_0, s37_1_1, s37_1_2, s37_1_3, s37_1_4, s37_1_5, s37_2_0, s37_2_1, s37_2_2, s37_2_3, s37_3_0, s37_3_1, s37_3_2, s37_4_0;
	wire s37_4_1, s37_5_0, s37_6_0, s37_7_0, s38_0_0, s38_0_1, s38_0_2, s38_0_3, s38_0_4, s38_0_5, s38_0_6, s38_0_7, s38_1_0, s38_1_1, s38_1_2, s38_1_3;
	wire s38_1_4, s38_1_5, s38_2_0, s38_2_1, s38_2_2, s38_2_3, s38_3_0, s38_3_1, s38_3_2, s38_4_0, s38_4_1, s38_5_0, s38_6_0, s38_7_0, s39_0_0, s39_0_1;
	wire s39_0_2, s39_0_3, s39_0_4, s39_0_5, s39_0_6, s39_0_7, s39_1_0, s39_1_1, s39_1_2, s39_1_3, s39_1_4, s39_2_0, s39_2_1, s39_2_2, s39_2_3, s39_3_0;
	wire s39_3_1, s39_3_2, s39_4_0, s39_4_1, s39_5_0, s39_6_0, s39_7_0, s3_0_0, s3_1_0, s3_2_0, s40_0_0, s40_0_1, s40_0_2, s40_0_3, s40_0_4, s40_0_5;
	wire s40_0_6, s40_0_7, s40_1_0, s40_1_1, s40_1_2, s40_1_3, s40_1_4, s40_2_0, s40_2_1, s40_2_2, s40_2_3, s40_3_0, s40_3_1, s40_3_2, s40_4_0, s40_4_1;
	wire s40_5_0, s40_6_0, s40_7_0, s41_0_0, s41_0_1, s41_0_2, s41_0_3, s41_0_4, s41_0_5, s41_0_6, s41_1_0, s41_1_1, s41_1_2, s41_1_3, s41_1_4, s41_2_0;
	wire s41_2_1, s41_2_2, s41_2_3, s41_3_0, s41_3_1, s41_3_2, s41_4_0, s41_4_1, s41_5_0, s41_6_0, s41_7_0, s42_0_0, s42_0_1, s42_0_2, s42_0_3, s42_0_4;
	wire s42_0_5, s42_0_6, s42_1_0, s42_1_1, s42_1_2, s42_1_3, s42_1_4, s42_2_0, s42_2_1, s42_2_2, s42_3_0, s42_3_1, s42_3_2, s42_4_0, s42_4_1, s42_5_0;
	wire s42_6_0, s42_7_0, s43_0_0, s43_0_1, s43_0_2, s43_0_3, s43_0_4, s43_0_5, s43_0_6, s43_1_0, s43_1_1, s43_1_2, s43_1_3, s43_1_4, s43_2_0, s43_2_1;
	wire s43_2_2, s43_3_0, s43_3_1, s43_4_0, s43_4_1, s43_5_0, s43_6_0, s43_7_0, s44_0_0, s44_0_1, s44_0_2, s44_0_3, s44_0_4, s44_0_5, s44_1_0, s44_1_1;
	wire s44_1_2, s44_1_3, s44_1_4, s44_2_0, s44_2_1, s44_2_2, s44_3_0, s44_3_1, s44_4_0, s44_4_1, s44_5_0, s44_6_0, s44_7_0, s45_0_0, s45_0_1, s45_0_2;
	wire s45_0_3, s45_0_4, s45_0_5, s45_1_0, s45_1_1, s45_1_2, s45_1_3, s45_2_0, s45_2_1, s45_2_2, s45_3_0, s45_3_1, s45_4_0, s45_5_0, s45_6_0, s45_7_0;
	wire s46_0_0, s46_0_1, s46_0_2, s46_0_3, s46_0_4, s46_0_5, s46_1_0, s46_1_1, s46_1_2, s46_1_3, s46_2_0, s46_2_1, s46_2_2, s46_3_0, s46_3_1, s46_4_0;
	wire s46_5_0, s46_6_0, s46_7_0, s47_0_0, s47_0_1, s47_0_2, s47_0_3, s47_0_4, s47_1_0, s47_1_1, s47_1_2, s47_1_3, s47_2_0, s47_2_1, s47_2_2, s47_3_0;
	wire s47_3_1, s47_4_0, s47_5_0, s47_6_0, s47_7_0, s48_0_0, s48_0_1, s48_0_2, s48_0_3, s48_0_4, s48_1_0, s48_1_1, s48_1_2, s48_2_0, s48_2_1, s48_2_2;
	wire s48_3_0, s48_3_1, s48_4_0, s48_5_0, s48_6_0, s48_7_0, s49_0_0, s49_0_1, s49_0_2, s49_0_3, s49_0_4, s49_1_0, s49_1_1, s49_1_2, s49_2_0, s49_2_1;
	wire s49_3_0, s49_3_1, s49_4_0, s49_5_0, s49_6_0, s49_7_0, s4_0_0, s4_0_1, s4_1_0, s4_2_0, s4_3_0, s50_0_0, s50_0_1, s50_0_2, s50_0_3, s50_1_0;
	wire s50_1_1, s50_1_2, s50_2_0, s50_2_1, s50_3_0, s50_3_1, s50_4_0, s50_5_0, s50_6_0, s50_7_0, s51_0_0, s51_0_1, s51_0_2, s51_0_3, s51_1_0, s51_1_1;
	wire s51_1_2, s51_2_0, s51_2_1, s51_3_0, s51_4_0, s51_5_0, s51_6_0, s51_7_0, s52_0_0, s52_0_1, s52_0_2, s52_0_3, s52_1_0, s52_1_1, s52_1_2, s52_2_0;
	wire s52_2_1, s52_3_0, s52_4_0, s52_5_0, s52_6_0, s52_7_0, s53_0_0, s53_0_1, s53_0_2, s53_1_0, s53_1_1, s53_1_2, s53_2_0, s53_2_1, s53_3_0, s53_4_0;
	wire s53_5_0, s53_6_0, s53_7_0, s54_0_0, s54_0_1, s54_0_2, s54_1_0, s54_1_1, s54_2_0, s54_2_1, s54_3_0, s54_4_0, s54_5_0, s54_6_0, s54_7_0, s55_0_0;
	wire s55_0_1, s55_0_2, s55_1_0, s55_1_1, s55_2_0, s55_3_0, s55_4_0, s55_5_0, s55_6_0, s55_7_0, s56_0_0, s56_0_1, s56_1_0, s56_1_1, s56_2_0, s56_3_0;
	wire s56_4_0, s56_5_0, s56_6_0, s56_7_0, s57_0_0, s57_0_1, s57_1_0, s57_2_0, s57_3_0, s57_4_0, s57_5_0, s57_6_0, s57_7_0, s58_0_0, s58_0_1, s58_1_0;
	wire s58_2_0, s58_3_0, s58_4_0, s58_5_0, s58_6_0, s58_7_0, s59_0_0, s59_1_0, s59_2_0, s59_3_0, s59_4_0, s59_5_0, s59_6_0, s59_7_0, s5_0_0, s5_0_1;
	wire s5_1_0, s5_2_0, s5_3_0, s5_4_0, s60_0_0, s60_1_0, s60_2_0, s60_3_0, s60_4_0, s60_5_0, s60_6_0, s60_7_0, s61_0_0, s61_1_0, s61_2_0, s61_3_0;
	wire s61_4_0, s61_5_0, s61_6_0, s61_7_0, s62_1_0, s62_2_0, s62_3_0, s62_4_0, s62_5_0, s62_6_0, s62_7_0, s63_2_0, s63_3_0, s63_4_0, s63_5_0, s63_6_0;
	wire s63_7_0, s6_0_0, s6_0_1, s6_1_0, s6_1_1, s6_2_0, s6_3_0, s6_4_0, s6_5_0, s7_0_0, s7_0_1, s7_0_2, s7_1_0, s7_1_1, s7_2_0, s7_3_0;
	wire s7_4_0, s7_5_0, s7_6_0, s8_0_0, s8_0_1, s8_0_2, s8_1_0, s8_1_1, s8_2_0, s8_3_0, s8_4_0, s8_5_0, s8_6_0, s8_7_0, s9_0_0, s9_0_1;
	wire s9_0_2, s9_1_0, s9_1_1, s9_2_0, s9_2_1, s9_3_0, s9_4_0, s9_5_0, s9_6_0, s9_7_0;
	
	wire cout, cout_a, cout_b;
	wire[63:0] x, y;
	wire[31:0] upperbits_a, upperbits_b, upperbits;
	wire xo_0, xo_1, xo_2, xo_3, xo_4, xo_5, xo_6, xo_7, xo_8, xo_9, xo_10, xo_11, xo_12, xo_13, xo_14, xo_15;
	wire o_0, o_1, o_2, o_3, o_4, n_0, xno_0, n_overflow;
	

	
	and and0_0(a0_0, B[0], A[0]);
	and and0_1(a0_1, B[0], A[1]);
	and and0_2(a0_2, B[0], A[2]);
	and and0_3(a0_3, B[0], A[3]);
	and and0_4(a0_4, B[0], A[4]);
	and and0_5(a0_5, B[0], A[5]);
	and and0_6(a0_6, B[0], A[6]);
	and and0_7(a0_7, B[0], A[7]);
	and and0_8(a0_8, B[0], A[8]);
	and and0_9(a0_9, B[0], A[9]);
	and and0_10(a0_10, B[0], A[10]);
	and and0_11(a0_11, B[0], A[11]);
	and and0_12(a0_12, B[0], A[12]);
	and and0_13(a0_13, B[0], A[13]);
	and and0_14(a0_14, B[0], A[14]);
	and and0_15(a0_15, B[0], A[15]);
	and and0_16(a0_16, B[0], A[16]);
	and and0_17(a0_17, B[0], A[17]);
	and and0_18(a0_18, B[0], A[18]);
	and and0_19(a0_19, B[0], A[19]);
	and and0_20(a0_20, B[0], A[20]);
	and and0_21(a0_21, B[0], A[21]);
	and and0_22(a0_22, B[0], A[22]);
	and and0_23(a0_23, B[0], A[23]);
	and and0_24(a0_24, B[0], A[24]);
	and and0_25(a0_25, B[0], A[25]);
	and and0_26(a0_26, B[0], A[26]);
	and and0_27(a0_27, B[0], A[27]);
	and and0_28(a0_28, B[0], A[28]);
	and and0_29(a0_29, B[0], A[29]);
	and and0_30(a0_30, B[0], A[30]);
	and and0_31(ap0_31, B[0], A[31]);
	and and1_1(a1_1, B[1], A[0]);
	and and1_2(a1_2, B[1], A[1]);
	and and1_3(a1_3, B[1], A[2]);
	and and1_4(a1_4, B[1], A[3]);
	and and1_5(a1_5, B[1], A[4]);
	and and1_6(a1_6, B[1], A[5]);
	and and1_7(a1_7, B[1], A[6]);
	and and1_8(a1_8, B[1], A[7]);
	and and1_9(a1_9, B[1], A[8]);
	and and1_10(a1_10, B[1], A[9]);
	and and1_11(a1_11, B[1], A[10]);
	and and1_12(a1_12, B[1], A[11]);
	and and1_13(a1_13, B[1], A[12]);
	and and1_14(a1_14, B[1], A[13]);
	and and1_15(a1_15, B[1], A[14]);
	and and1_16(a1_16, B[1], A[15]);
	and and1_17(a1_17, B[1], A[16]);
	and and1_18(a1_18, B[1], A[17]);
	and and1_19(a1_19, B[1], A[18]);
	and and1_20(a1_20, B[1], A[19]);
	and and1_21(a1_21, B[1], A[20]);
	and and1_22(a1_22, B[1], A[21]);
	and and1_23(a1_23, B[1], A[22]);
	and and1_24(a1_24, B[1], A[23]);
	and and1_25(a1_25, B[1], A[24]);
	and and1_26(a1_26, B[1], A[25]);
	and and1_27(a1_27, B[1], A[26]);
	and and1_28(a1_28, B[1], A[27]);
	and and1_29(a1_29, B[1], A[28]);
	and and1_30(a1_30, B[1], A[29]);
	and and1_31(a1_31, B[1], A[30]);
	and and1_32(ap1_32, B[1], A[31]);
	and and2_2(a2_2, B[2], A[0]);
	and and2_3(a2_3, B[2], A[1]);
	and and2_4(a2_4, B[2], A[2]);
	and and2_5(a2_5, B[2], A[3]);
	and and2_6(a2_6, B[2], A[4]);
	and and2_7(a2_7, B[2], A[5]);
	and and2_8(a2_8, B[2], A[6]);
	and and2_9(a2_9, B[2], A[7]);
	and and2_10(a2_10, B[2], A[8]);
	and and2_11(a2_11, B[2], A[9]);
	and and2_12(a2_12, B[2], A[10]);
	and and2_13(a2_13, B[2], A[11]);
	and and2_14(a2_14, B[2], A[12]);
	and and2_15(a2_15, B[2], A[13]);
	and and2_16(a2_16, B[2], A[14]);
	and and2_17(a2_17, B[2], A[15]);
	and and2_18(a2_18, B[2], A[16]);
	and and2_19(a2_19, B[2], A[17]);
	and and2_20(a2_20, B[2], A[18]);
	and and2_21(a2_21, B[2], A[19]);
	and and2_22(a2_22, B[2], A[20]);
	and and2_23(a2_23, B[2], A[21]);
	and and2_24(a2_24, B[2], A[22]);
	and and2_25(a2_25, B[2], A[23]);
	and and2_26(a2_26, B[2], A[24]);
	and and2_27(a2_27, B[2], A[25]);
	and and2_28(a2_28, B[2], A[26]);
	and and2_29(a2_29, B[2], A[27]);
	and and2_30(a2_30, B[2], A[28]);
	and and2_31(a2_31, B[2], A[29]);
	and and2_32(a2_32, B[2], A[30]);
	and and2_33(ap2_33, B[2], A[31]);
	and and3_3(a3_3, B[3], A[0]);
	and and3_4(a3_4, B[3], A[1]);
	and and3_5(a3_5, B[3], A[2]);
	and and3_6(a3_6, B[3], A[3]);
	and and3_7(a3_7, B[3], A[4]);
	and and3_8(a3_8, B[3], A[5]);
	and and3_9(a3_9, B[3], A[6]);
	and and3_10(a3_10, B[3], A[7]);
	and and3_11(a3_11, B[3], A[8]);
	and and3_12(a3_12, B[3], A[9]);
	and and3_13(a3_13, B[3], A[10]);
	and and3_14(a3_14, B[3], A[11]);
	and and3_15(a3_15, B[3], A[12]);
	and and3_16(a3_16, B[3], A[13]);
	and and3_17(a3_17, B[3], A[14]);
	and and3_18(a3_18, B[3], A[15]);
	and and3_19(a3_19, B[3], A[16]);
	and and3_20(a3_20, B[3], A[17]);
	and and3_21(a3_21, B[3], A[18]);
	and and3_22(a3_22, B[3], A[19]);
	and and3_23(a3_23, B[3], A[20]);
	and and3_24(a3_24, B[3], A[21]);
	and and3_25(a3_25, B[3], A[22]);
	and and3_26(a3_26, B[3], A[23]);
	and and3_27(a3_27, B[3], A[24]);
	and and3_28(a3_28, B[3], A[25]);
	and and3_29(a3_29, B[3], A[26]);
	and and3_30(a3_30, B[3], A[27]);
	and and3_31(a3_31, B[3], A[28]);
	and and3_32(a3_32, B[3], A[29]);
	and and3_33(a3_33, B[3], A[30]);
	and and3_34(ap3_34, B[3], A[31]);
	and and4_4(a4_4, B[4], A[0]);
	and and4_5(a4_5, B[4], A[1]);
	and and4_6(a4_6, B[4], A[2]);
	and and4_7(a4_7, B[4], A[3]);
	and and4_8(a4_8, B[4], A[4]);
	and and4_9(a4_9, B[4], A[5]);
	and and4_10(a4_10, B[4], A[6]);
	and and4_11(a4_11, B[4], A[7]);
	and and4_12(a4_12, B[4], A[8]);
	and and4_13(a4_13, B[4], A[9]);
	and and4_14(a4_14, B[4], A[10]);
	and and4_15(a4_15, B[4], A[11]);
	and and4_16(a4_16, B[4], A[12]);
	and and4_17(a4_17, B[4], A[13]);
	and and4_18(a4_18, B[4], A[14]);
	and and4_19(a4_19, B[4], A[15]);
	and and4_20(a4_20, B[4], A[16]);
	and and4_21(a4_21, B[4], A[17]);
	and and4_22(a4_22, B[4], A[18]);
	and and4_23(a4_23, B[4], A[19]);
	and and4_24(a4_24, B[4], A[20]);
	and and4_25(a4_25, B[4], A[21]);
	and and4_26(a4_26, B[4], A[22]);
	and and4_27(a4_27, B[4], A[23]);
	and and4_28(a4_28, B[4], A[24]);
	and and4_29(a4_29, B[4], A[25]);
	and and4_30(a4_30, B[4], A[26]);
	and and4_31(a4_31, B[4], A[27]);
	and and4_32(a4_32, B[4], A[28]);
	and and4_33(a4_33, B[4], A[29]);
	and and4_34(a4_34, B[4], A[30]);
	and and4_35(ap4_35, B[4], A[31]);
	and and5_5(a5_5, B[5], A[0]);
	and and5_6(a5_6, B[5], A[1]);
	and and5_7(a5_7, B[5], A[2]);
	and and5_8(a5_8, B[5], A[3]);
	and and5_9(a5_9, B[5], A[4]);
	and and5_10(a5_10, B[5], A[5]);
	and and5_11(a5_11, B[5], A[6]);
	and and5_12(a5_12, B[5], A[7]);
	and and5_13(a5_13, B[5], A[8]);
	and and5_14(a5_14, B[5], A[9]);
	and and5_15(a5_15, B[5], A[10]);
	and and5_16(a5_16, B[5], A[11]);
	and and5_17(a5_17, B[5], A[12]);
	and and5_18(a5_18, B[5], A[13]);
	and and5_19(a5_19, B[5], A[14]);
	and and5_20(a5_20, B[5], A[15]);
	and and5_21(a5_21, B[5], A[16]);
	and and5_22(a5_22, B[5], A[17]);
	and and5_23(a5_23, B[5], A[18]);
	and and5_24(a5_24, B[5], A[19]);
	and and5_25(a5_25, B[5], A[20]);
	and and5_26(a5_26, B[5], A[21]);
	and and5_27(a5_27, B[5], A[22]);
	and and5_28(a5_28, B[5], A[23]);
	and and5_29(a5_29, B[5], A[24]);
	and and5_30(a5_30, B[5], A[25]);
	and and5_31(a5_31, B[5], A[26]);
	and and5_32(a5_32, B[5], A[27]);
	and and5_33(a5_33, B[5], A[28]);
	and and5_34(a5_34, B[5], A[29]);
	and and5_35(a5_35, B[5], A[30]);
	and and5_36(ap5_36, B[5], A[31]);
	and and6_6(a6_6, B[6], A[0]);
	and and6_7(a6_7, B[6], A[1]);
	and and6_8(a6_8, B[6], A[2]);
	and and6_9(a6_9, B[6], A[3]);
	and and6_10(a6_10, B[6], A[4]);
	and and6_11(a6_11, B[6], A[5]);
	and and6_12(a6_12, B[6], A[6]);
	and and6_13(a6_13, B[6], A[7]);
	and and6_14(a6_14, B[6], A[8]);
	and and6_15(a6_15, B[6], A[9]);
	and and6_16(a6_16, B[6], A[10]);
	and and6_17(a6_17, B[6], A[11]);
	and and6_18(a6_18, B[6], A[12]);
	and and6_19(a6_19, B[6], A[13]);
	and and6_20(a6_20, B[6], A[14]);
	and and6_21(a6_21, B[6], A[15]);
	and and6_22(a6_22, B[6], A[16]);
	and and6_23(a6_23, B[6], A[17]);
	and and6_24(a6_24, B[6], A[18]);
	and and6_25(a6_25, B[6], A[19]);
	and and6_26(a6_26, B[6], A[20]);
	and and6_27(a6_27, B[6], A[21]);
	and and6_28(a6_28, B[6], A[22]);
	and and6_29(a6_29, B[6], A[23]);
	and and6_30(a6_30, B[6], A[24]);
	and and6_31(a6_31, B[6], A[25]);
	and and6_32(a6_32, B[6], A[26]);
	and and6_33(a6_33, B[6], A[27]);
	and and6_34(a6_34, B[6], A[28]);
	and and6_35(a6_35, B[6], A[29]);
	and and6_36(a6_36, B[6], A[30]);
	and and6_37(ap6_37, B[6], A[31]);
	and and7_7(a7_7, B[7], A[0]);
	and and7_8(a7_8, B[7], A[1]);
	and and7_9(a7_9, B[7], A[2]);
	and and7_10(a7_10, B[7], A[3]);
	and and7_11(a7_11, B[7], A[4]);
	and and7_12(a7_12, B[7], A[5]);
	and and7_13(a7_13, B[7], A[6]);
	and and7_14(a7_14, B[7], A[7]);
	and and7_15(a7_15, B[7], A[8]);
	and and7_16(a7_16, B[7], A[9]);
	and and7_17(a7_17, B[7], A[10]);
	and and7_18(a7_18, B[7], A[11]);
	and and7_19(a7_19, B[7], A[12]);
	and and7_20(a7_20, B[7], A[13]);
	and and7_21(a7_21, B[7], A[14]);
	and and7_22(a7_22, B[7], A[15]);
	and and7_23(a7_23, B[7], A[16]);
	and and7_24(a7_24, B[7], A[17]);
	and and7_25(a7_25, B[7], A[18]);
	and and7_26(a7_26, B[7], A[19]);
	and and7_27(a7_27, B[7], A[20]);
	and and7_28(a7_28, B[7], A[21]);
	and and7_29(a7_29, B[7], A[22]);
	and and7_30(a7_30, B[7], A[23]);
	and and7_31(a7_31, B[7], A[24]);
	and and7_32(a7_32, B[7], A[25]);
	and and7_33(a7_33, B[7], A[26]);
	and and7_34(a7_34, B[7], A[27]);
	and and7_35(a7_35, B[7], A[28]);
	and and7_36(a7_36, B[7], A[29]);
	and and7_37(a7_37, B[7], A[30]);
	and and7_38(ap7_38, B[7], A[31]);
	and and8_8(a8_8, B[8], A[0]);
	and and8_9(a8_9, B[8], A[1]);
	and and8_10(a8_10, B[8], A[2]);
	and and8_11(a8_11, B[8], A[3]);
	and and8_12(a8_12, B[8], A[4]);
	and and8_13(a8_13, B[8], A[5]);
	and and8_14(a8_14, B[8], A[6]);
	and and8_15(a8_15, B[8], A[7]);
	and and8_16(a8_16, B[8], A[8]);
	and and8_17(a8_17, B[8], A[9]);
	and and8_18(a8_18, B[8], A[10]);
	and and8_19(a8_19, B[8], A[11]);
	and and8_20(a8_20, B[8], A[12]);
	and and8_21(a8_21, B[8], A[13]);
	and and8_22(a8_22, B[8], A[14]);
	and and8_23(a8_23, B[8], A[15]);
	and and8_24(a8_24, B[8], A[16]);
	and and8_25(a8_25, B[8], A[17]);
	and and8_26(a8_26, B[8], A[18]);
	and and8_27(a8_27, B[8], A[19]);
	and and8_28(a8_28, B[8], A[20]);
	and and8_29(a8_29, B[8], A[21]);
	and and8_30(a8_30, B[8], A[22]);
	and and8_31(a8_31, B[8], A[23]);
	and and8_32(a8_32, B[8], A[24]);
	and and8_33(a8_33, B[8], A[25]);
	and and8_34(a8_34, B[8], A[26]);
	and and8_35(a8_35, B[8], A[27]);
	and and8_36(a8_36, B[8], A[28]);
	and and8_37(a8_37, B[8], A[29]);
	and and8_38(a8_38, B[8], A[30]);
	and and8_39(ap8_39, B[8], A[31]);
	and and9_9(a9_9, B[9], A[0]);
	and and9_10(a9_10, B[9], A[1]);
	and and9_11(a9_11, B[9], A[2]);
	and and9_12(a9_12, B[9], A[3]);
	and and9_13(a9_13, B[9], A[4]);
	and and9_14(a9_14, B[9], A[5]);
	and and9_15(a9_15, B[9], A[6]);
	and and9_16(a9_16, B[9], A[7]);
	and and9_17(a9_17, B[9], A[8]);
	and and9_18(a9_18, B[9], A[9]);
	and and9_19(a9_19, B[9], A[10]);
	and and9_20(a9_20, B[9], A[11]);
	and and9_21(a9_21, B[9], A[12]);
	and and9_22(a9_22, B[9], A[13]);
	and and9_23(a9_23, B[9], A[14]);
	and and9_24(a9_24, B[9], A[15]);
	and and9_25(a9_25, B[9], A[16]);
	and and9_26(a9_26, B[9], A[17]);
	and and9_27(a9_27, B[9], A[18]);
	and and9_28(a9_28, B[9], A[19]);
	and and9_29(a9_29, B[9], A[20]);
	and and9_30(a9_30, B[9], A[21]);
	and and9_31(a9_31, B[9], A[22]);
	and and9_32(a9_32, B[9], A[23]);
	and and9_33(a9_33, B[9], A[24]);
	and and9_34(a9_34, B[9], A[25]);
	and and9_35(a9_35, B[9], A[26]);
	and and9_36(a9_36, B[9], A[27]);
	and and9_37(a9_37, B[9], A[28]);
	and and9_38(a9_38, B[9], A[29]);
	and and9_39(a9_39, B[9], A[30]);
	and and9_40(ap9_40, B[9], A[31]);
	and and10_10(a10_10, B[10], A[0]);
	and and10_11(a10_11, B[10], A[1]);
	and and10_12(a10_12, B[10], A[2]);
	and and10_13(a10_13, B[10], A[3]);
	and and10_14(a10_14, B[10], A[4]);
	and and10_15(a10_15, B[10], A[5]);
	and and10_16(a10_16, B[10], A[6]);
	and and10_17(a10_17, B[10], A[7]);
	and and10_18(a10_18, B[10], A[8]);
	and and10_19(a10_19, B[10], A[9]);
	and and10_20(a10_20, B[10], A[10]);
	and and10_21(a10_21, B[10], A[11]);
	and and10_22(a10_22, B[10], A[12]);
	and and10_23(a10_23, B[10], A[13]);
	and and10_24(a10_24, B[10], A[14]);
	and and10_25(a10_25, B[10], A[15]);
	and and10_26(a10_26, B[10], A[16]);
	and and10_27(a10_27, B[10], A[17]);
	and and10_28(a10_28, B[10], A[18]);
	and and10_29(a10_29, B[10], A[19]);
	and and10_30(a10_30, B[10], A[20]);
	and and10_31(a10_31, B[10], A[21]);
	and and10_32(a10_32, B[10], A[22]);
	and and10_33(a10_33, B[10], A[23]);
	and and10_34(a10_34, B[10], A[24]);
	and and10_35(a10_35, B[10], A[25]);
	and and10_36(a10_36, B[10], A[26]);
	and and10_37(a10_37, B[10], A[27]);
	and and10_38(a10_38, B[10], A[28]);
	and and10_39(a10_39, B[10], A[29]);
	and and10_40(a10_40, B[10], A[30]);
	and and10_41(ap10_41, B[10], A[31]);
	and and11_11(a11_11, B[11], A[0]);
	and and11_12(a11_12, B[11], A[1]);
	and and11_13(a11_13, B[11], A[2]);
	and and11_14(a11_14, B[11], A[3]);
	and and11_15(a11_15, B[11], A[4]);
	and and11_16(a11_16, B[11], A[5]);
	and and11_17(a11_17, B[11], A[6]);
	and and11_18(a11_18, B[11], A[7]);
	and and11_19(a11_19, B[11], A[8]);
	and and11_20(a11_20, B[11], A[9]);
	and and11_21(a11_21, B[11], A[10]);
	and and11_22(a11_22, B[11], A[11]);
	and and11_23(a11_23, B[11], A[12]);
	and and11_24(a11_24, B[11], A[13]);
	and and11_25(a11_25, B[11], A[14]);
	and and11_26(a11_26, B[11], A[15]);
	and and11_27(a11_27, B[11], A[16]);
	and and11_28(a11_28, B[11], A[17]);
	and and11_29(a11_29, B[11], A[18]);
	and and11_30(a11_30, B[11], A[19]);
	and and11_31(a11_31, B[11], A[20]);
	and and11_32(a11_32, B[11], A[21]);
	and and11_33(a11_33, B[11], A[22]);
	and and11_34(a11_34, B[11], A[23]);
	and and11_35(a11_35, B[11], A[24]);
	and and11_36(a11_36, B[11], A[25]);
	and and11_37(a11_37, B[11], A[26]);
	and and11_38(a11_38, B[11], A[27]);
	and and11_39(a11_39, B[11], A[28]);
	and and11_40(a11_40, B[11], A[29]);
	and and11_41(a11_41, B[11], A[30]);
	and and11_42(ap11_42, B[11], A[31]);
	and and12_12(a12_12, B[12], A[0]);
	and and12_13(a12_13, B[12], A[1]);
	and and12_14(a12_14, B[12], A[2]);
	and and12_15(a12_15, B[12], A[3]);
	and and12_16(a12_16, B[12], A[4]);
	and and12_17(a12_17, B[12], A[5]);
	and and12_18(a12_18, B[12], A[6]);
	and and12_19(a12_19, B[12], A[7]);
	and and12_20(a12_20, B[12], A[8]);
	and and12_21(a12_21, B[12], A[9]);
	and and12_22(a12_22, B[12], A[10]);
	and and12_23(a12_23, B[12], A[11]);
	and and12_24(a12_24, B[12], A[12]);
	and and12_25(a12_25, B[12], A[13]);
	and and12_26(a12_26, B[12], A[14]);
	and and12_27(a12_27, B[12], A[15]);
	and and12_28(a12_28, B[12], A[16]);
	and and12_29(a12_29, B[12], A[17]);
	and and12_30(a12_30, B[12], A[18]);
	and and12_31(a12_31, B[12], A[19]);
	and and12_32(a12_32, B[12], A[20]);
	and and12_33(a12_33, B[12], A[21]);
	and and12_34(a12_34, B[12], A[22]);
	and and12_35(a12_35, B[12], A[23]);
	and and12_36(a12_36, B[12], A[24]);
	and and12_37(a12_37, B[12], A[25]);
	and and12_38(a12_38, B[12], A[26]);
	and and12_39(a12_39, B[12], A[27]);
	and and12_40(a12_40, B[12], A[28]);
	and and12_41(a12_41, B[12], A[29]);
	and and12_42(a12_42, B[12], A[30]);
	and and12_43(ap12_43, B[12], A[31]);
	and and13_13(a13_13, B[13], A[0]);
	and and13_14(a13_14, B[13], A[1]);
	and and13_15(a13_15, B[13], A[2]);
	and and13_16(a13_16, B[13], A[3]);
	and and13_17(a13_17, B[13], A[4]);
	and and13_18(a13_18, B[13], A[5]);
	and and13_19(a13_19, B[13], A[6]);
	and and13_20(a13_20, B[13], A[7]);
	and and13_21(a13_21, B[13], A[8]);
	and and13_22(a13_22, B[13], A[9]);
	and and13_23(a13_23, B[13], A[10]);
	and and13_24(a13_24, B[13], A[11]);
	and and13_25(a13_25, B[13], A[12]);
	and and13_26(a13_26, B[13], A[13]);
	and and13_27(a13_27, B[13], A[14]);
	and and13_28(a13_28, B[13], A[15]);
	and and13_29(a13_29, B[13], A[16]);
	and and13_30(a13_30, B[13], A[17]);
	and and13_31(a13_31, B[13], A[18]);
	and and13_32(a13_32, B[13], A[19]);
	and and13_33(a13_33, B[13], A[20]);
	and and13_34(a13_34, B[13], A[21]);
	and and13_35(a13_35, B[13], A[22]);
	and and13_36(a13_36, B[13], A[23]);
	and and13_37(a13_37, B[13], A[24]);
	and and13_38(a13_38, B[13], A[25]);
	and and13_39(a13_39, B[13], A[26]);
	and and13_40(a13_40, B[13], A[27]);
	and and13_41(a13_41, B[13], A[28]);
	and and13_42(a13_42, B[13], A[29]);
	and and13_43(a13_43, B[13], A[30]);
	and and13_44(ap13_44, B[13], A[31]);
	and and14_14(a14_14, B[14], A[0]);
	and and14_15(a14_15, B[14], A[1]);
	and and14_16(a14_16, B[14], A[2]);
	and and14_17(a14_17, B[14], A[3]);
	and and14_18(a14_18, B[14], A[4]);
	and and14_19(a14_19, B[14], A[5]);
	and and14_20(a14_20, B[14], A[6]);
	and and14_21(a14_21, B[14], A[7]);
	and and14_22(a14_22, B[14], A[8]);
	and and14_23(a14_23, B[14], A[9]);
	and and14_24(a14_24, B[14], A[10]);
	and and14_25(a14_25, B[14], A[11]);
	and and14_26(a14_26, B[14], A[12]);
	and and14_27(a14_27, B[14], A[13]);
	and and14_28(a14_28, B[14], A[14]);
	and and14_29(a14_29, B[14], A[15]);
	and and14_30(a14_30, B[14], A[16]);
	and and14_31(a14_31, B[14], A[17]);
	and and14_32(a14_32, B[14], A[18]);
	and and14_33(a14_33, B[14], A[19]);
	and and14_34(a14_34, B[14], A[20]);
	and and14_35(a14_35, B[14], A[21]);
	and and14_36(a14_36, B[14], A[22]);
	and and14_37(a14_37, B[14], A[23]);
	and and14_38(a14_38, B[14], A[24]);
	and and14_39(a14_39, B[14], A[25]);
	and and14_40(a14_40, B[14], A[26]);
	and and14_41(a14_41, B[14], A[27]);
	and and14_42(a14_42, B[14], A[28]);
	and and14_43(a14_43, B[14], A[29]);
	and and14_44(a14_44, B[14], A[30]);
	and and14_45(ap14_45, B[14], A[31]);
	and and15_15(a15_15, B[15], A[0]);
	and and15_16(a15_16, B[15], A[1]);
	and and15_17(a15_17, B[15], A[2]);
	and and15_18(a15_18, B[15], A[3]);
	and and15_19(a15_19, B[15], A[4]);
	and and15_20(a15_20, B[15], A[5]);
	and and15_21(a15_21, B[15], A[6]);
	and and15_22(a15_22, B[15], A[7]);
	and and15_23(a15_23, B[15], A[8]);
	and and15_24(a15_24, B[15], A[9]);
	and and15_25(a15_25, B[15], A[10]);
	and and15_26(a15_26, B[15], A[11]);
	and and15_27(a15_27, B[15], A[12]);
	and and15_28(a15_28, B[15], A[13]);
	and and15_29(a15_29, B[15], A[14]);
	and and15_30(a15_30, B[15], A[15]);
	and and15_31(a15_31, B[15], A[16]);
	and and15_32(a15_32, B[15], A[17]);
	and and15_33(a15_33, B[15], A[18]);
	and and15_34(a15_34, B[15], A[19]);
	and and15_35(a15_35, B[15], A[20]);
	and and15_36(a15_36, B[15], A[21]);
	and and15_37(a15_37, B[15], A[22]);
	and and15_38(a15_38, B[15], A[23]);
	and and15_39(a15_39, B[15], A[24]);
	and and15_40(a15_40, B[15], A[25]);
	and and15_41(a15_41, B[15], A[26]);
	and and15_42(a15_42, B[15], A[27]);
	and and15_43(a15_43, B[15], A[28]);
	and and15_44(a15_44, B[15], A[29]);
	and and15_45(a15_45, B[15], A[30]);
	and and15_46(ap15_46, B[15], A[31]);
	and and16_16(a16_16, B[16], A[0]);
	and and16_17(a16_17, B[16], A[1]);
	and and16_18(a16_18, B[16], A[2]);
	and and16_19(a16_19, B[16], A[3]);
	and and16_20(a16_20, B[16], A[4]);
	and and16_21(a16_21, B[16], A[5]);
	and and16_22(a16_22, B[16], A[6]);
	and and16_23(a16_23, B[16], A[7]);
	and and16_24(a16_24, B[16], A[8]);
	and and16_25(a16_25, B[16], A[9]);
	and and16_26(a16_26, B[16], A[10]);
	and and16_27(a16_27, B[16], A[11]);
	and and16_28(a16_28, B[16], A[12]);
	and and16_29(a16_29, B[16], A[13]);
	and and16_30(a16_30, B[16], A[14]);
	and and16_31(a16_31, B[16], A[15]);
	and and16_32(a16_32, B[16], A[16]);
	and and16_33(a16_33, B[16], A[17]);
	and and16_34(a16_34, B[16], A[18]);
	and and16_35(a16_35, B[16], A[19]);
	and and16_36(a16_36, B[16], A[20]);
	and and16_37(a16_37, B[16], A[21]);
	and and16_38(a16_38, B[16], A[22]);
	and and16_39(a16_39, B[16], A[23]);
	and and16_40(a16_40, B[16], A[24]);
	and and16_41(a16_41, B[16], A[25]);
	and and16_42(a16_42, B[16], A[26]);
	and and16_43(a16_43, B[16], A[27]);
	and and16_44(a16_44, B[16], A[28]);
	and and16_45(a16_45, B[16], A[29]);
	and and16_46(a16_46, B[16], A[30]);
	and and16_47(ap16_47, B[16], A[31]);
	and and17_17(a17_17, B[17], A[0]);
	and and17_18(a17_18, B[17], A[1]);
	and and17_19(a17_19, B[17], A[2]);
	and and17_20(a17_20, B[17], A[3]);
	and and17_21(a17_21, B[17], A[4]);
	and and17_22(a17_22, B[17], A[5]);
	and and17_23(a17_23, B[17], A[6]);
	and and17_24(a17_24, B[17], A[7]);
	and and17_25(a17_25, B[17], A[8]);
	and and17_26(a17_26, B[17], A[9]);
	and and17_27(a17_27, B[17], A[10]);
	and and17_28(a17_28, B[17], A[11]);
	and and17_29(a17_29, B[17], A[12]);
	and and17_30(a17_30, B[17], A[13]);
	and and17_31(a17_31, B[17], A[14]);
	and and17_32(a17_32, B[17], A[15]);
	and and17_33(a17_33, B[17], A[16]);
	and and17_34(a17_34, B[17], A[17]);
	and and17_35(a17_35, B[17], A[18]);
	and and17_36(a17_36, B[17], A[19]);
	and and17_37(a17_37, B[17], A[20]);
	and and17_38(a17_38, B[17], A[21]);
	and and17_39(a17_39, B[17], A[22]);
	and and17_40(a17_40, B[17], A[23]);
	and and17_41(a17_41, B[17], A[24]);
	and and17_42(a17_42, B[17], A[25]);
	and and17_43(a17_43, B[17], A[26]);
	and and17_44(a17_44, B[17], A[27]);
	and and17_45(a17_45, B[17], A[28]);
	and and17_46(a17_46, B[17], A[29]);
	and and17_47(a17_47, B[17], A[30]);
	and and17_48(ap17_48, B[17], A[31]);
	and and18_18(a18_18, B[18], A[0]);
	and and18_19(a18_19, B[18], A[1]);
	and and18_20(a18_20, B[18], A[2]);
	and and18_21(a18_21, B[18], A[3]);
	and and18_22(a18_22, B[18], A[4]);
	and and18_23(a18_23, B[18], A[5]);
	and and18_24(a18_24, B[18], A[6]);
	and and18_25(a18_25, B[18], A[7]);
	and and18_26(a18_26, B[18], A[8]);
	and and18_27(a18_27, B[18], A[9]);
	and and18_28(a18_28, B[18], A[10]);
	and and18_29(a18_29, B[18], A[11]);
	and and18_30(a18_30, B[18], A[12]);
	and and18_31(a18_31, B[18], A[13]);
	and and18_32(a18_32, B[18], A[14]);
	and and18_33(a18_33, B[18], A[15]);
	and and18_34(a18_34, B[18], A[16]);
	and and18_35(a18_35, B[18], A[17]);
	and and18_36(a18_36, B[18], A[18]);
	and and18_37(a18_37, B[18], A[19]);
	and and18_38(a18_38, B[18], A[20]);
	and and18_39(a18_39, B[18], A[21]);
	and and18_40(a18_40, B[18], A[22]);
	and and18_41(a18_41, B[18], A[23]);
	and and18_42(a18_42, B[18], A[24]);
	and and18_43(a18_43, B[18], A[25]);
	and and18_44(a18_44, B[18], A[26]);
	and and18_45(a18_45, B[18], A[27]);
	and and18_46(a18_46, B[18], A[28]);
	and and18_47(a18_47, B[18], A[29]);
	and and18_48(a18_48, B[18], A[30]);
	and and18_49(ap18_49, B[18], A[31]);
	and and19_19(a19_19, B[19], A[0]);
	and and19_20(a19_20, B[19], A[1]);
	and and19_21(a19_21, B[19], A[2]);
	and and19_22(a19_22, B[19], A[3]);
	and and19_23(a19_23, B[19], A[4]);
	and and19_24(a19_24, B[19], A[5]);
	and and19_25(a19_25, B[19], A[6]);
	and and19_26(a19_26, B[19], A[7]);
	and and19_27(a19_27, B[19], A[8]);
	and and19_28(a19_28, B[19], A[9]);
	and and19_29(a19_29, B[19], A[10]);
	and and19_30(a19_30, B[19], A[11]);
	and and19_31(a19_31, B[19], A[12]);
	and and19_32(a19_32, B[19], A[13]);
	and and19_33(a19_33, B[19], A[14]);
	and and19_34(a19_34, B[19], A[15]);
	and and19_35(a19_35, B[19], A[16]);
	and and19_36(a19_36, B[19], A[17]);
	and and19_37(a19_37, B[19], A[18]);
	and and19_38(a19_38, B[19], A[19]);
	and and19_39(a19_39, B[19], A[20]);
	and and19_40(a19_40, B[19], A[21]);
	and and19_41(a19_41, B[19], A[22]);
	and and19_42(a19_42, B[19], A[23]);
	and and19_43(a19_43, B[19], A[24]);
	and and19_44(a19_44, B[19], A[25]);
	and and19_45(a19_45, B[19], A[26]);
	and and19_46(a19_46, B[19], A[27]);
	and and19_47(a19_47, B[19], A[28]);
	and and19_48(a19_48, B[19], A[29]);
	and and19_49(a19_49, B[19], A[30]);
	and and19_50(ap19_50, B[19], A[31]);
	and and20_20(a20_20, B[20], A[0]);
	and and20_21(a20_21, B[20], A[1]);
	and and20_22(a20_22, B[20], A[2]);
	and and20_23(a20_23, B[20], A[3]);
	and and20_24(a20_24, B[20], A[4]);
	and and20_25(a20_25, B[20], A[5]);
	and and20_26(a20_26, B[20], A[6]);
	and and20_27(a20_27, B[20], A[7]);
	and and20_28(a20_28, B[20], A[8]);
	and and20_29(a20_29, B[20], A[9]);
	and and20_30(a20_30, B[20], A[10]);
	and and20_31(a20_31, B[20], A[11]);
	and and20_32(a20_32, B[20], A[12]);
	and and20_33(a20_33, B[20], A[13]);
	and and20_34(a20_34, B[20], A[14]);
	and and20_35(a20_35, B[20], A[15]);
	and and20_36(a20_36, B[20], A[16]);
	and and20_37(a20_37, B[20], A[17]);
	and and20_38(a20_38, B[20], A[18]);
	and and20_39(a20_39, B[20], A[19]);
	and and20_40(a20_40, B[20], A[20]);
	and and20_41(a20_41, B[20], A[21]);
	and and20_42(a20_42, B[20], A[22]);
	and and20_43(a20_43, B[20], A[23]);
	and and20_44(a20_44, B[20], A[24]);
	and and20_45(a20_45, B[20], A[25]);
	and and20_46(a20_46, B[20], A[26]);
	and and20_47(a20_47, B[20], A[27]);
	and and20_48(a20_48, B[20], A[28]);
	and and20_49(a20_49, B[20], A[29]);
	and and20_50(a20_50, B[20], A[30]);
	and and20_51(ap20_51, B[20], A[31]);
	and and21_21(a21_21, B[21], A[0]);
	and and21_22(a21_22, B[21], A[1]);
	and and21_23(a21_23, B[21], A[2]);
	and and21_24(a21_24, B[21], A[3]);
	and and21_25(a21_25, B[21], A[4]);
	and and21_26(a21_26, B[21], A[5]);
	and and21_27(a21_27, B[21], A[6]);
	and and21_28(a21_28, B[21], A[7]);
	and and21_29(a21_29, B[21], A[8]);
	and and21_30(a21_30, B[21], A[9]);
	and and21_31(a21_31, B[21], A[10]);
	and and21_32(a21_32, B[21], A[11]);
	and and21_33(a21_33, B[21], A[12]);
	and and21_34(a21_34, B[21], A[13]);
	and and21_35(a21_35, B[21], A[14]);
	and and21_36(a21_36, B[21], A[15]);
	and and21_37(a21_37, B[21], A[16]);
	and and21_38(a21_38, B[21], A[17]);
	and and21_39(a21_39, B[21], A[18]);
	and and21_40(a21_40, B[21], A[19]);
	and and21_41(a21_41, B[21], A[20]);
	and and21_42(a21_42, B[21], A[21]);
	and and21_43(a21_43, B[21], A[22]);
	and and21_44(a21_44, B[21], A[23]);
	and and21_45(a21_45, B[21], A[24]);
	and and21_46(a21_46, B[21], A[25]);
	and and21_47(a21_47, B[21], A[26]);
	and and21_48(a21_48, B[21], A[27]);
	and and21_49(a21_49, B[21], A[28]);
	and and21_50(a21_50, B[21], A[29]);
	and and21_51(a21_51, B[21], A[30]);
	and and21_52(ap21_52, B[21], A[31]);
	and and22_22(a22_22, B[22], A[0]);
	and and22_23(a22_23, B[22], A[1]);
	and and22_24(a22_24, B[22], A[2]);
	and and22_25(a22_25, B[22], A[3]);
	and and22_26(a22_26, B[22], A[4]);
	and and22_27(a22_27, B[22], A[5]);
	and and22_28(a22_28, B[22], A[6]);
	and and22_29(a22_29, B[22], A[7]);
	and and22_30(a22_30, B[22], A[8]);
	and and22_31(a22_31, B[22], A[9]);
	and and22_32(a22_32, B[22], A[10]);
	and and22_33(a22_33, B[22], A[11]);
	and and22_34(a22_34, B[22], A[12]);
	and and22_35(a22_35, B[22], A[13]);
	and and22_36(a22_36, B[22], A[14]);
	and and22_37(a22_37, B[22], A[15]);
	and and22_38(a22_38, B[22], A[16]);
	and and22_39(a22_39, B[22], A[17]);
	and and22_40(a22_40, B[22], A[18]);
	and and22_41(a22_41, B[22], A[19]);
	and and22_42(a22_42, B[22], A[20]);
	and and22_43(a22_43, B[22], A[21]);
	and and22_44(a22_44, B[22], A[22]);
	and and22_45(a22_45, B[22], A[23]);
	and and22_46(a22_46, B[22], A[24]);
	and and22_47(a22_47, B[22], A[25]);
	and and22_48(a22_48, B[22], A[26]);
	and and22_49(a22_49, B[22], A[27]);
	and and22_50(a22_50, B[22], A[28]);
	and and22_51(a22_51, B[22], A[29]);
	and and22_52(a22_52, B[22], A[30]);
	and and22_53(ap22_53, B[22], A[31]);
	and and23_23(a23_23, B[23], A[0]);
	and and23_24(a23_24, B[23], A[1]);
	and and23_25(a23_25, B[23], A[2]);
	and and23_26(a23_26, B[23], A[3]);
	and and23_27(a23_27, B[23], A[4]);
	and and23_28(a23_28, B[23], A[5]);
	and and23_29(a23_29, B[23], A[6]);
	and and23_30(a23_30, B[23], A[7]);
	and and23_31(a23_31, B[23], A[8]);
	and and23_32(a23_32, B[23], A[9]);
	and and23_33(a23_33, B[23], A[10]);
	and and23_34(a23_34, B[23], A[11]);
	and and23_35(a23_35, B[23], A[12]);
	and and23_36(a23_36, B[23], A[13]);
	and and23_37(a23_37, B[23], A[14]);
	and and23_38(a23_38, B[23], A[15]);
	and and23_39(a23_39, B[23], A[16]);
	and and23_40(a23_40, B[23], A[17]);
	and and23_41(a23_41, B[23], A[18]);
	and and23_42(a23_42, B[23], A[19]);
	and and23_43(a23_43, B[23], A[20]);
	and and23_44(a23_44, B[23], A[21]);
	and and23_45(a23_45, B[23], A[22]);
	and and23_46(a23_46, B[23], A[23]);
	and and23_47(a23_47, B[23], A[24]);
	and and23_48(a23_48, B[23], A[25]);
	and and23_49(a23_49, B[23], A[26]);
	and and23_50(a23_50, B[23], A[27]);
	and and23_51(a23_51, B[23], A[28]);
	and and23_52(a23_52, B[23], A[29]);
	and and23_53(a23_53, B[23], A[30]);
	and and23_54(ap23_54, B[23], A[31]);
	and and24_24(a24_24, B[24], A[0]);
	and and24_25(a24_25, B[24], A[1]);
	and and24_26(a24_26, B[24], A[2]);
	and and24_27(a24_27, B[24], A[3]);
	and and24_28(a24_28, B[24], A[4]);
	and and24_29(a24_29, B[24], A[5]);
	and and24_30(a24_30, B[24], A[6]);
	and and24_31(a24_31, B[24], A[7]);
	and and24_32(a24_32, B[24], A[8]);
	and and24_33(a24_33, B[24], A[9]);
	and and24_34(a24_34, B[24], A[10]);
	and and24_35(a24_35, B[24], A[11]);
	and and24_36(a24_36, B[24], A[12]);
	and and24_37(a24_37, B[24], A[13]);
	and and24_38(a24_38, B[24], A[14]);
	and and24_39(a24_39, B[24], A[15]);
	and and24_40(a24_40, B[24], A[16]);
	and and24_41(a24_41, B[24], A[17]);
	and and24_42(a24_42, B[24], A[18]);
	and and24_43(a24_43, B[24], A[19]);
	and and24_44(a24_44, B[24], A[20]);
	and and24_45(a24_45, B[24], A[21]);
	and and24_46(a24_46, B[24], A[22]);
	and and24_47(a24_47, B[24], A[23]);
	and and24_48(a24_48, B[24], A[24]);
	and and24_49(a24_49, B[24], A[25]);
	and and24_50(a24_50, B[24], A[26]);
	and and24_51(a24_51, B[24], A[27]);
	and and24_52(a24_52, B[24], A[28]);
	and and24_53(a24_53, B[24], A[29]);
	and and24_54(a24_54, B[24], A[30]);
	and and24_55(ap24_55, B[24], A[31]);
	and and25_25(a25_25, B[25], A[0]);
	and and25_26(a25_26, B[25], A[1]);
	and and25_27(a25_27, B[25], A[2]);
	and and25_28(a25_28, B[25], A[3]);
	and and25_29(a25_29, B[25], A[4]);
	and and25_30(a25_30, B[25], A[5]);
	and and25_31(a25_31, B[25], A[6]);
	and and25_32(a25_32, B[25], A[7]);
	and and25_33(a25_33, B[25], A[8]);
	and and25_34(a25_34, B[25], A[9]);
	and and25_35(a25_35, B[25], A[10]);
	and and25_36(a25_36, B[25], A[11]);
	and and25_37(a25_37, B[25], A[12]);
	and and25_38(a25_38, B[25], A[13]);
	and and25_39(a25_39, B[25], A[14]);
	and and25_40(a25_40, B[25], A[15]);
	and and25_41(a25_41, B[25], A[16]);
	and and25_42(a25_42, B[25], A[17]);
	and and25_43(a25_43, B[25], A[18]);
	and and25_44(a25_44, B[25], A[19]);
	and and25_45(a25_45, B[25], A[20]);
	and and25_46(a25_46, B[25], A[21]);
	and and25_47(a25_47, B[25], A[22]);
	and and25_48(a25_48, B[25], A[23]);
	and and25_49(a25_49, B[25], A[24]);
	and and25_50(a25_50, B[25], A[25]);
	and and25_51(a25_51, B[25], A[26]);
	and and25_52(a25_52, B[25], A[27]);
	and and25_53(a25_53, B[25], A[28]);
	and and25_54(a25_54, B[25], A[29]);
	and and25_55(a25_55, B[25], A[30]);
	and and25_56(ap25_56, B[25], A[31]);
	and and26_26(a26_26, B[26], A[0]);
	and and26_27(a26_27, B[26], A[1]);
	and and26_28(a26_28, B[26], A[2]);
	and and26_29(a26_29, B[26], A[3]);
	and and26_30(a26_30, B[26], A[4]);
	and and26_31(a26_31, B[26], A[5]);
	and and26_32(a26_32, B[26], A[6]);
	and and26_33(a26_33, B[26], A[7]);
	and and26_34(a26_34, B[26], A[8]);
	and and26_35(a26_35, B[26], A[9]);
	and and26_36(a26_36, B[26], A[10]);
	and and26_37(a26_37, B[26], A[11]);
	and and26_38(a26_38, B[26], A[12]);
	and and26_39(a26_39, B[26], A[13]);
	and and26_40(a26_40, B[26], A[14]);
	and and26_41(a26_41, B[26], A[15]);
	and and26_42(a26_42, B[26], A[16]);
	and and26_43(a26_43, B[26], A[17]);
	and and26_44(a26_44, B[26], A[18]);
	and and26_45(a26_45, B[26], A[19]);
	and and26_46(a26_46, B[26], A[20]);
	and and26_47(a26_47, B[26], A[21]);
	and and26_48(a26_48, B[26], A[22]);
	and and26_49(a26_49, B[26], A[23]);
	and and26_50(a26_50, B[26], A[24]);
	and and26_51(a26_51, B[26], A[25]);
	and and26_52(a26_52, B[26], A[26]);
	and and26_53(a26_53, B[26], A[27]);
	and and26_54(a26_54, B[26], A[28]);
	and and26_55(a26_55, B[26], A[29]);
	and and26_56(a26_56, B[26], A[30]);
	and and26_57(ap26_57, B[26], A[31]);
	and and27_27(a27_27, B[27], A[0]);
	and and27_28(a27_28, B[27], A[1]);
	and and27_29(a27_29, B[27], A[2]);
	and and27_30(a27_30, B[27], A[3]);
	and and27_31(a27_31, B[27], A[4]);
	and and27_32(a27_32, B[27], A[5]);
	and and27_33(a27_33, B[27], A[6]);
	and and27_34(a27_34, B[27], A[7]);
	and and27_35(a27_35, B[27], A[8]);
	and and27_36(a27_36, B[27], A[9]);
	and and27_37(a27_37, B[27], A[10]);
	and and27_38(a27_38, B[27], A[11]);
	and and27_39(a27_39, B[27], A[12]);
	and and27_40(a27_40, B[27], A[13]);
	and and27_41(a27_41, B[27], A[14]);
	and and27_42(a27_42, B[27], A[15]);
	and and27_43(a27_43, B[27], A[16]);
	and and27_44(a27_44, B[27], A[17]);
	and and27_45(a27_45, B[27], A[18]);
	and and27_46(a27_46, B[27], A[19]);
	and and27_47(a27_47, B[27], A[20]);
	and and27_48(a27_48, B[27], A[21]);
	and and27_49(a27_49, B[27], A[22]);
	and and27_50(a27_50, B[27], A[23]);
	and and27_51(a27_51, B[27], A[24]);
	and and27_52(a27_52, B[27], A[25]);
	and and27_53(a27_53, B[27], A[26]);
	and and27_54(a27_54, B[27], A[27]);
	and and27_55(a27_55, B[27], A[28]);
	and and27_56(a27_56, B[27], A[29]);
	and and27_57(a27_57, B[27], A[30]);
	and and27_58(ap27_58, B[27], A[31]);
	and and28_28(a28_28, B[28], A[0]);
	and and28_29(a28_29, B[28], A[1]);
	and and28_30(a28_30, B[28], A[2]);
	and and28_31(a28_31, B[28], A[3]);
	and and28_32(a28_32, B[28], A[4]);
	and and28_33(a28_33, B[28], A[5]);
	and and28_34(a28_34, B[28], A[6]);
	and and28_35(a28_35, B[28], A[7]);
	and and28_36(a28_36, B[28], A[8]);
	and and28_37(a28_37, B[28], A[9]);
	and and28_38(a28_38, B[28], A[10]);
	and and28_39(a28_39, B[28], A[11]);
	and and28_40(a28_40, B[28], A[12]);
	and and28_41(a28_41, B[28], A[13]);
	and and28_42(a28_42, B[28], A[14]);
	and and28_43(a28_43, B[28], A[15]);
	and and28_44(a28_44, B[28], A[16]);
	and and28_45(a28_45, B[28], A[17]);
	and and28_46(a28_46, B[28], A[18]);
	and and28_47(a28_47, B[28], A[19]);
	and and28_48(a28_48, B[28], A[20]);
	and and28_49(a28_49, B[28], A[21]);
	and and28_50(a28_50, B[28], A[22]);
	and and28_51(a28_51, B[28], A[23]);
	and and28_52(a28_52, B[28], A[24]);
	and and28_53(a28_53, B[28], A[25]);
	and and28_54(a28_54, B[28], A[26]);
	and and28_55(a28_55, B[28], A[27]);
	and and28_56(a28_56, B[28], A[28]);
	and and28_57(a28_57, B[28], A[29]);
	and and28_58(a28_58, B[28], A[30]);
	and and28_59(ap28_59, B[28], A[31]);
	and and29_29(a29_29, B[29], A[0]);
	and and29_30(a29_30, B[29], A[1]);
	and and29_31(a29_31, B[29], A[2]);
	and and29_32(a29_32, B[29], A[3]);
	and and29_33(a29_33, B[29], A[4]);
	and and29_34(a29_34, B[29], A[5]);
	and and29_35(a29_35, B[29], A[6]);
	and and29_36(a29_36, B[29], A[7]);
	and and29_37(a29_37, B[29], A[8]);
	and and29_38(a29_38, B[29], A[9]);
	and and29_39(a29_39, B[29], A[10]);
	and and29_40(a29_40, B[29], A[11]);
	and and29_41(a29_41, B[29], A[12]);
	and and29_42(a29_42, B[29], A[13]);
	and and29_43(a29_43, B[29], A[14]);
	and and29_44(a29_44, B[29], A[15]);
	and and29_45(a29_45, B[29], A[16]);
	and and29_46(a29_46, B[29], A[17]);
	and and29_47(a29_47, B[29], A[18]);
	and and29_48(a29_48, B[29], A[19]);
	and and29_49(a29_49, B[29], A[20]);
	and and29_50(a29_50, B[29], A[21]);
	and and29_51(a29_51, B[29], A[22]);
	and and29_52(a29_52, B[29], A[23]);
	and and29_53(a29_53, B[29], A[24]);
	and and29_54(a29_54, B[29], A[25]);
	and and29_55(a29_55, B[29], A[26]);
	and and29_56(a29_56, B[29], A[27]);
	and and29_57(a29_57, B[29], A[28]);
	and and29_58(a29_58, B[29], A[29]);
	and and29_59(a29_59, B[29], A[30]);
	and and29_60(ap29_60, B[29], A[31]);
	and and30_30(a30_30, B[30], A[0]);
	and and30_31(a30_31, B[30], A[1]);
	and and30_32(a30_32, B[30], A[2]);
	and and30_33(a30_33, B[30], A[3]);
	and and30_34(a30_34, B[30], A[4]);
	and and30_35(a30_35, B[30], A[5]);
	and and30_36(a30_36, B[30], A[6]);
	and and30_37(a30_37, B[30], A[7]);
	and and30_38(a30_38, B[30], A[8]);
	and and30_39(a30_39, B[30], A[9]);
	and and30_40(a30_40, B[30], A[10]);
	and and30_41(a30_41, B[30], A[11]);
	and and30_42(a30_42, B[30], A[12]);
	and and30_43(a30_43, B[30], A[13]);
	and and30_44(a30_44, B[30], A[14]);
	and and30_45(a30_45, B[30], A[15]);
	and and30_46(a30_46, B[30], A[16]);
	and and30_47(a30_47, B[30], A[17]);
	and and30_48(a30_48, B[30], A[18]);
	and and30_49(a30_49, B[30], A[19]);
	and and30_50(a30_50, B[30], A[20]);
	and and30_51(a30_51, B[30], A[21]);
	and and30_52(a30_52, B[30], A[22]);
	and and30_53(a30_53, B[30], A[23]);
	and and30_54(a30_54, B[30], A[24]);
	and and30_55(a30_55, B[30], A[25]);
	and and30_56(a30_56, B[30], A[26]);
	and and30_57(a30_57, B[30], A[27]);
	and and30_58(a30_58, B[30], A[28]);
	and and30_59(a30_59, B[30], A[29]);
	and and30_60(a30_60, B[30], A[30]);
	and and30_61(ap30_61, B[30], A[31]);
	and and31_31(ap31_31, B[31], A[0]);
	and and31_32(ap31_32, B[31], A[1]);
	and and31_33(ap31_33, B[31], A[2]);
	and and31_34(ap31_34, B[31], A[3]);
	and and31_35(ap31_35, B[31], A[4]);
	and and31_36(ap31_36, B[31], A[5]);
	and and31_37(ap31_37, B[31], A[6]);
	and and31_38(ap31_38, B[31], A[7]);
	and and31_39(ap31_39, B[31], A[8]);
	and and31_40(ap31_40, B[31], A[9]);
	and and31_41(ap31_41, B[31], A[10]);
	and and31_42(ap31_42, B[31], A[11]);
	and and31_43(ap31_43, B[31], A[12]);
	and and31_44(ap31_44, B[31], A[13]);
	and and31_45(ap31_45, B[31], A[14]);
	and and31_46(ap31_46, B[31], A[15]);
	and and31_47(ap31_47, B[31], A[16]);
	and and31_48(ap31_48, B[31], A[17]);
	and and31_49(ap31_49, B[31], A[18]);
	and and31_50(ap31_50, B[31], A[19]);
	and and31_51(ap31_51, B[31], A[20]);
	and and31_52(ap31_52, B[31], A[21]);
	and and31_53(ap31_53, B[31], A[22]);
	and and31_54(ap31_54, B[31], A[23]);
	and and31_55(ap31_55, B[31], A[24]);
	and and31_56(ap31_56, B[31], A[25]);
	and and31_57(ap31_57, B[31], A[26]);
	and and31_58(ap31_58, B[31], A[27]);
	and and31_59(ap31_59, B[31], A[28]);
	and and31_60(ap31_60, B[31], A[29]);
	and and31_61(ap31_61, B[31], A[30]);
	and and31_62(a31_62, B[31], A[31]);

	not not0_31(a0_31, ap0_31);
	not not1_32(a1_32, ap1_32);
	not not2_33(a2_33, ap2_33);
	not not3_34(a3_34, ap3_34);
	not not4_35(a4_35, ap4_35);
	not not5_36(a5_36, ap5_36);
	not not6_37(a6_37, ap6_37);
	not not7_38(a7_38, ap7_38);
	not not8_39(a8_39, ap8_39);
	not not9_40(a9_40, ap9_40);
	not not10_41(a10_41, ap10_41);
	not not11_42(a11_42, ap11_42);
	not not12_43(a12_43, ap12_43);
	not not13_44(a13_44, ap13_44);
	not not14_45(a14_45, ap14_45);
	not not15_46(a15_46, ap15_46);
	not not16_47(a16_47, ap16_47);
	not not17_48(a17_48, ap17_48);
	not not18_49(a18_49, ap18_49);
	not not19_50(a19_50, ap19_50);
	not not20_51(a20_51, ap20_51);
	not not21_52(a21_52, ap21_52);
	not not22_53(a22_53, ap22_53);
	not not23_54(a23_54, ap23_54);
	not not24_55(a24_55, ap24_55);
	not not25_56(a25_56, ap25_56);
	not not26_57(a26_57, ap26_57);
	not not27_58(a27_58, ap27_58);
	not not28_59(a28_59, ap28_59);
	not not29_60(a29_60, ap29_60);
	not not30_61(a30_61, ap30_61);
	not not31_31(a31_31, ap31_31);
	not not31_32(a31_32, ap31_32);
	not not31_33(a31_33, ap31_33);
	not not31_34(a31_34, ap31_34);
	not not31_35(a31_35, ap31_35);
	not not31_36(a31_36, ap31_36);
	not not31_37(a31_37, ap31_37);
	not not31_38(a31_38, ap31_38);
	not not31_39(a31_39, ap31_39);
	not not31_40(a31_40, ap31_40);
	not not31_41(a31_41, ap31_41);
	not not31_42(a31_42, ap31_42);
	not not31_43(a31_43, ap31_43);
	not not31_44(a31_44, ap31_44);
	not not31_45(a31_45, ap31_45);
	not not31_46(a31_46, ap31_46);
	not not31_47(a31_47, ap31_47);
	not not31_48(a31_48, ap31_48);
	not not31_49(a31_49, ap31_49);
	not not31_50(a31_50, ap31_50);
	not not31_51(a31_51, ap31_51);
	not not31_52(a31_52, ap31_52);
	not not31_53(a31_53, ap31_53);
	not not31_54(a31_54, ap31_54);
	not not31_55(a31_55, ap31_55);
	not not31_56(a31_56, ap31_56);
	not not31_57(a31_57, ap31_57);
	not not31_58(a31_58, ap31_58);
	not not31_59(a31_59, ap31_59);
	not not31_60(a31_60, ap31_60);
	not not31_61(a31_61, ap31_61);

	half_adder ha1_0_0(a0_1, a1_1, s1_0_0, c1_0_0);
	full_adder ad2_0_0(a0_2, a1_2, a2_2, s2_0_0, c2_0_0);
	full_adder ad3_0_0(a0_3, a1_3, a2_3, s3_0_0, c3_0_0);
	full_adder ad4_0_0(a0_4, a1_4, a2_4, s4_0_0, c4_0_0);
	half_adder ha4_0_1(a3_4, a4_4, s4_0_1, c4_0_1);
	full_adder ad5_0_0(a0_5, a1_5, a2_5, s5_0_0, c5_0_0);
	full_adder ad5_0_1(a3_5, a4_5, a5_5, s5_0_1, c5_0_1);
	full_adder ad6_0_0(a0_6, a1_6, a2_6, s6_0_0, c6_0_0);
	full_adder ad6_0_1(a3_6, a4_6, a5_6, s6_0_1, c6_0_1);
	full_adder ad7_0_0(a0_7, a1_7, a2_7, s7_0_0, c7_0_0);
	full_adder ad7_0_1(a3_7, a4_7, a5_7, s7_0_1, c7_0_1);
	half_adder ha7_0_2(a6_7, a7_7, s7_0_2, c7_0_2);
	full_adder ad8_0_0(a0_8, a1_8, a2_8, s8_0_0, c8_0_0);
	full_adder ad8_0_1(a3_8, a4_8, a5_8, s8_0_1, c8_0_1);
	full_adder ad8_0_2(a6_8, a7_8, a8_8, s8_0_2, c8_0_2);
	full_adder ad9_0_0(a0_9, a1_9, a2_9, s9_0_0, c9_0_0);
	full_adder ad9_0_1(a3_9, a4_9, a5_9, s9_0_1, c9_0_1);
	full_adder ad9_0_2(a6_9, a7_9, a8_9, s9_0_2, c9_0_2);
	full_adder ad10_0_0(a0_10, a1_10, a2_10, s10_0_0, c10_0_0);
	full_adder ad10_0_1(a3_10, a4_10, a5_10, s10_0_1, c10_0_1);
	full_adder ad10_0_2(a6_10, a7_10, a8_10, s10_0_2, c10_0_2);
	half_adder ha10_0_3(a9_10, a10_10, s10_0_3, c10_0_3);
	full_adder ad11_0_0(a0_11, a1_11, a2_11, s11_0_0, c11_0_0);
	full_adder ad11_0_1(a3_11, a4_11, a5_11, s11_0_1, c11_0_1);
	full_adder ad11_0_2(a6_11, a7_11, a8_11, s11_0_2, c11_0_2);
	full_adder ad11_0_3(a9_11, a10_11, a11_11, s11_0_3, c11_0_3);
	full_adder ad12_0_0(a0_12, a1_12, a2_12, s12_0_0, c12_0_0);
	full_adder ad12_0_1(a3_12, a4_12, a5_12, s12_0_1, c12_0_1);
	full_adder ad12_0_2(a6_12, a7_12, a8_12, s12_0_2, c12_0_2);
	full_adder ad12_0_3(a9_12, a10_12, a11_12, s12_0_3, c12_0_3);
	full_adder ad13_0_0(a0_13, a1_13, a2_13, s13_0_0, c13_0_0);
	full_adder ad13_0_1(a3_13, a4_13, a5_13, s13_0_1, c13_0_1);
	full_adder ad13_0_2(a6_13, a7_13, a8_13, s13_0_2, c13_0_2);
	full_adder ad13_0_3(a9_13, a10_13, a11_13, s13_0_3, c13_0_3);
	half_adder ha13_0_4(a12_13, a13_13, s13_0_4, c13_0_4);
	full_adder ad14_0_0(a0_14, a1_14, a2_14, s14_0_0, c14_0_0);
	full_adder ad14_0_1(a3_14, a4_14, a5_14, s14_0_1, c14_0_1);
	full_adder ad14_0_2(a6_14, a7_14, a8_14, s14_0_2, c14_0_2);
	full_adder ad14_0_3(a9_14, a10_14, a11_14, s14_0_3, c14_0_3);
	full_adder ad14_0_4(a12_14, a13_14, a14_14, s14_0_4, c14_0_4);
	full_adder ad15_0_0(a0_15, a1_15, a2_15, s15_0_0, c15_0_0);
	full_adder ad15_0_1(a3_15, a4_15, a5_15, s15_0_1, c15_0_1);
	full_adder ad15_0_2(a6_15, a7_15, a8_15, s15_0_2, c15_0_2);
	full_adder ad15_0_3(a9_15, a10_15, a11_15, s15_0_3, c15_0_3);
	full_adder ad15_0_4(a12_15, a13_15, a14_15, s15_0_4, c15_0_4);
	full_adder ad16_0_0(a0_16, a1_16, a2_16, s16_0_0, c16_0_0);
	full_adder ad16_0_1(a3_16, a4_16, a5_16, s16_0_1, c16_0_1);
	full_adder ad16_0_2(a6_16, a7_16, a8_16, s16_0_2, c16_0_2);
	full_adder ad16_0_3(a9_16, a10_16, a11_16, s16_0_3, c16_0_3);
	full_adder ad16_0_4(a12_16, a13_16, a14_16, s16_0_4, c16_0_4);
	half_adder ha16_0_5(a15_16, a16_16, s16_0_5, c16_0_5);
	full_adder ad17_0_0(a0_17, a1_17, a2_17, s17_0_0, c17_0_0);
	full_adder ad17_0_1(a3_17, a4_17, a5_17, s17_0_1, c17_0_1);
	full_adder ad17_0_2(a6_17, a7_17, a8_17, s17_0_2, c17_0_2);
	full_adder ad17_0_3(a9_17, a10_17, a11_17, s17_0_3, c17_0_3);
	full_adder ad17_0_4(a12_17, a13_17, a14_17, s17_0_4, c17_0_4);
	full_adder ad17_0_5(a15_17, a16_17, a17_17, s17_0_5, c17_0_5);
	full_adder ad18_0_0(a0_18, a1_18, a2_18, s18_0_0, c18_0_0);
	full_adder ad18_0_1(a3_18, a4_18, a5_18, s18_0_1, c18_0_1);
	full_adder ad18_0_2(a6_18, a7_18, a8_18, s18_0_2, c18_0_2);
	full_adder ad18_0_3(a9_18, a10_18, a11_18, s18_0_3, c18_0_3);
	full_adder ad18_0_4(a12_18, a13_18, a14_18, s18_0_4, c18_0_4);
	full_adder ad18_0_5(a15_18, a16_18, a17_18, s18_0_5, c18_0_5);
	full_adder ad19_0_0(a0_19, a1_19, a2_19, s19_0_0, c19_0_0);
	full_adder ad19_0_1(a3_19, a4_19, a5_19, s19_0_1, c19_0_1);
	full_adder ad19_0_2(a6_19, a7_19, a8_19, s19_0_2, c19_0_2);
	full_adder ad19_0_3(a9_19, a10_19, a11_19, s19_0_3, c19_0_3);
	full_adder ad19_0_4(a12_19, a13_19, a14_19, s19_0_4, c19_0_4);
	full_adder ad19_0_5(a15_19, a16_19, a17_19, s19_0_5, c19_0_5);
	half_adder ha19_0_6(a18_19, a19_19, s19_0_6, c19_0_6);
	full_adder ad20_0_0(a0_20, a1_20, a2_20, s20_0_0, c20_0_0);
	full_adder ad20_0_1(a3_20, a4_20, a5_20, s20_0_1, c20_0_1);
	full_adder ad20_0_2(a6_20, a7_20, a8_20, s20_0_2, c20_0_2);
	full_adder ad20_0_3(a9_20, a10_20, a11_20, s20_0_3, c20_0_3);
	full_adder ad20_0_4(a12_20, a13_20, a14_20, s20_0_4, c20_0_4);
	full_adder ad20_0_5(a15_20, a16_20, a17_20, s20_0_5, c20_0_5);
	full_adder ad20_0_6(a18_20, a19_20, a20_20, s20_0_6, c20_0_6);
	full_adder ad21_0_0(a0_21, a1_21, a2_21, s21_0_0, c21_0_0);
	full_adder ad21_0_1(a3_21, a4_21, a5_21, s21_0_1, c21_0_1);
	full_adder ad21_0_2(a6_21, a7_21, a8_21, s21_0_2, c21_0_2);
	full_adder ad21_0_3(a9_21, a10_21, a11_21, s21_0_3, c21_0_3);
	full_adder ad21_0_4(a12_21, a13_21, a14_21, s21_0_4, c21_0_4);
	full_adder ad21_0_5(a15_21, a16_21, a17_21, s21_0_5, c21_0_5);
	full_adder ad21_0_6(a18_21, a19_21, a20_21, s21_0_6, c21_0_6);
	full_adder ad22_0_0(a0_22, a1_22, a2_22, s22_0_0, c22_0_0);
	full_adder ad22_0_1(a3_22, a4_22, a5_22, s22_0_1, c22_0_1);
	full_adder ad22_0_2(a6_22, a7_22, a8_22, s22_0_2, c22_0_2);
	full_adder ad22_0_3(a9_22, a10_22, a11_22, s22_0_3, c22_0_3);
	full_adder ad22_0_4(a12_22, a13_22, a14_22, s22_0_4, c22_0_4);
	full_adder ad22_0_5(a15_22, a16_22, a17_22, s22_0_5, c22_0_5);
	full_adder ad22_0_6(a18_22, a19_22, a20_22, s22_0_6, c22_0_6);
	half_adder ha22_0_7(a21_22, a22_22, s22_0_7, c22_0_7);
	full_adder ad23_0_0(a0_23, a1_23, a2_23, s23_0_0, c23_0_0);
	full_adder ad23_0_1(a3_23, a4_23, a5_23, s23_0_1, c23_0_1);
	full_adder ad23_0_2(a6_23, a7_23, a8_23, s23_0_2, c23_0_2);
	full_adder ad23_0_3(a9_23, a10_23, a11_23, s23_0_3, c23_0_3);
	full_adder ad23_0_4(a12_23, a13_23, a14_23, s23_0_4, c23_0_4);
	full_adder ad23_0_5(a15_23, a16_23, a17_23, s23_0_5, c23_0_5);
	full_adder ad23_0_6(a18_23, a19_23, a20_23, s23_0_6, c23_0_6);
	full_adder ad23_0_7(a21_23, a22_23, a23_23, s23_0_7, c23_0_7);
	full_adder ad24_0_0(a0_24, a1_24, a2_24, s24_0_0, c24_0_0);
	full_adder ad24_0_1(a3_24, a4_24, a5_24, s24_0_1, c24_0_1);
	full_adder ad24_0_2(a6_24, a7_24, a8_24, s24_0_2, c24_0_2);
	full_adder ad24_0_3(a9_24, a10_24, a11_24, s24_0_3, c24_0_3);
	full_adder ad24_0_4(a12_24, a13_24, a14_24, s24_0_4, c24_0_4);
	full_adder ad24_0_5(a15_24, a16_24, a17_24, s24_0_5, c24_0_5);
	full_adder ad24_0_6(a18_24, a19_24, a20_24, s24_0_6, c24_0_6);
	full_adder ad24_0_7(a21_24, a22_24, a23_24, s24_0_7, c24_0_7);
	full_adder ad25_0_0(a0_25, a1_25, a2_25, s25_0_0, c25_0_0);
	full_adder ad25_0_1(a3_25, a4_25, a5_25, s25_0_1, c25_0_1);
	full_adder ad25_0_2(a6_25, a7_25, a8_25, s25_0_2, c25_0_2);
	full_adder ad25_0_3(a9_25, a10_25, a11_25, s25_0_3, c25_0_3);
	full_adder ad25_0_4(a12_25, a13_25, a14_25, s25_0_4, c25_0_4);
	full_adder ad25_0_5(a15_25, a16_25, a17_25, s25_0_5, c25_0_5);
	full_adder ad25_0_6(a18_25, a19_25, a20_25, s25_0_6, c25_0_6);
	full_adder ad25_0_7(a21_25, a22_25, a23_25, s25_0_7, c25_0_7);
	half_adder ha25_0_8(a24_25, a25_25, s25_0_8, c25_0_8);
	full_adder ad26_0_0(a0_26, a1_26, a2_26, s26_0_0, c26_0_0);
	full_adder ad26_0_1(a3_26, a4_26, a5_26, s26_0_1, c26_0_1);
	full_adder ad26_0_2(a6_26, a7_26, a8_26, s26_0_2, c26_0_2);
	full_adder ad26_0_3(a9_26, a10_26, a11_26, s26_0_3, c26_0_3);
	full_adder ad26_0_4(a12_26, a13_26, a14_26, s26_0_4, c26_0_4);
	full_adder ad26_0_5(a15_26, a16_26, a17_26, s26_0_5, c26_0_5);
	full_adder ad26_0_6(a18_26, a19_26, a20_26, s26_0_6, c26_0_6);
	full_adder ad26_0_7(a21_26, a22_26, a23_26, s26_0_7, c26_0_7);
	full_adder ad26_0_8(a24_26, a25_26, a26_26, s26_0_8, c26_0_8);
	full_adder ad27_0_0(a0_27, a1_27, a2_27, s27_0_0, c27_0_0);
	full_adder ad27_0_1(a3_27, a4_27, a5_27, s27_0_1, c27_0_1);
	full_adder ad27_0_2(a6_27, a7_27, a8_27, s27_0_2, c27_0_2);
	full_adder ad27_0_3(a9_27, a10_27, a11_27, s27_0_3, c27_0_3);
	full_adder ad27_0_4(a12_27, a13_27, a14_27, s27_0_4, c27_0_4);
	full_adder ad27_0_5(a15_27, a16_27, a17_27, s27_0_5, c27_0_5);
	full_adder ad27_0_6(a18_27, a19_27, a20_27, s27_0_6, c27_0_6);
	full_adder ad27_0_7(a21_27, a22_27, a23_27, s27_0_7, c27_0_7);
	full_adder ad27_0_8(a24_27, a25_27, a26_27, s27_0_8, c27_0_8);
	full_adder ad28_0_0(a0_28, a1_28, a2_28, s28_0_0, c28_0_0);
	full_adder ad28_0_1(a3_28, a4_28, a5_28, s28_0_1, c28_0_1);
	full_adder ad28_0_2(a6_28, a7_28, a8_28, s28_0_2, c28_0_2);
	full_adder ad28_0_3(a9_28, a10_28, a11_28, s28_0_3, c28_0_3);
	full_adder ad28_0_4(a12_28, a13_28, a14_28, s28_0_4, c28_0_4);
	full_adder ad28_0_5(a15_28, a16_28, a17_28, s28_0_5, c28_0_5);
	full_adder ad28_0_6(a18_28, a19_28, a20_28, s28_0_6, c28_0_6);
	full_adder ad28_0_7(a21_28, a22_28, a23_28, s28_0_7, c28_0_7);
	full_adder ad28_0_8(a24_28, a25_28, a26_28, s28_0_8, c28_0_8);
	half_adder ha28_0_9(a27_28, a28_28, s28_0_9, c28_0_9);
	full_adder ad29_0_0(a0_29, a1_29, a2_29, s29_0_0, c29_0_0);
	full_adder ad29_0_1(a3_29, a4_29, a5_29, s29_0_1, c29_0_1);
	full_adder ad29_0_2(a6_29, a7_29, a8_29, s29_0_2, c29_0_2);
	full_adder ad29_0_3(a9_29, a10_29, a11_29, s29_0_3, c29_0_3);
	full_adder ad29_0_4(a12_29, a13_29, a14_29, s29_0_4, c29_0_4);
	full_adder ad29_0_5(a15_29, a16_29, a17_29, s29_0_5, c29_0_5);
	full_adder ad29_0_6(a18_29, a19_29, a20_29, s29_0_6, c29_0_6);
	full_adder ad29_0_7(a21_29, a22_29, a23_29, s29_0_7, c29_0_7);
	full_adder ad29_0_8(a24_29, a25_29, a26_29, s29_0_8, c29_0_8);
	full_adder ad29_0_9(a27_29, a28_29, a29_29, s29_0_9, c29_0_9);
	full_adder ad30_0_0(a0_30, a1_30, a2_30, s30_0_0, c30_0_0);
	full_adder ad30_0_1(a3_30, a4_30, a5_30, s30_0_1, c30_0_1);
	full_adder ad30_0_2(a6_30, a7_30, a8_30, s30_0_2, c30_0_2);
	full_adder ad30_0_3(a9_30, a10_30, a11_30, s30_0_3, c30_0_3);
	full_adder ad30_0_4(a12_30, a13_30, a14_30, s30_0_4, c30_0_4);
	full_adder ad30_0_5(a15_30, a16_30, a17_30, s30_0_5, c30_0_5);
	full_adder ad30_0_6(a18_30, a19_30, a20_30, s30_0_6, c30_0_6);
	full_adder ad30_0_7(a21_30, a22_30, a23_30, s30_0_7, c30_0_7);
	full_adder ad30_0_8(a24_30, a25_30, a26_30, s30_0_8, c30_0_8);
	full_adder ad30_0_9(a27_30, a28_30, a29_30, s30_0_9, c30_0_9);
	full_adder ad31_0_0(a0_31, a1_31, a2_31, s31_0_0, c31_0_0);
	full_adder ad31_0_1(a3_31, a4_31, a5_31, s31_0_1, c31_0_1);
	full_adder ad31_0_2(a6_31, a7_31, a8_31, s31_0_2, c31_0_2);
	full_adder ad31_0_3(a9_31, a10_31, a11_31, s31_0_3, c31_0_3);
	full_adder ad31_0_4(a12_31, a13_31, a14_31, s31_0_4, c31_0_4);
	full_adder ad31_0_5(a15_31, a16_31, a17_31, s31_0_5, c31_0_5);
	full_adder ad31_0_6(a18_31, a19_31, a20_31, s31_0_6, c31_0_6);
	full_adder ad31_0_7(a21_31, a22_31, a23_31, s31_0_7, c31_0_7);
	full_adder ad31_0_8(a24_31, a25_31, a26_31, s31_0_8, c31_0_8);
	full_adder ad31_0_9(a27_31, a28_31, a29_31, s31_0_9, c31_0_9);
	half_adder ha31_0_10(a30_31, a31_31, s31_0_10, c31_0_10);
	full_adder ad32_0_0(1'b1, a1_32, a2_32, s32_0_0, c32_0_0);
	full_adder ad32_0_1(a3_32, a4_32, a5_32, s32_0_1, c32_0_1);
	full_adder ad32_0_2(a6_32, a7_32, a8_32, s32_0_2, c32_0_2);
	full_adder ad32_0_3(a9_32, a10_32, a11_32, s32_0_3, c32_0_3);
	full_adder ad32_0_4(a12_32, a13_32, a14_32, s32_0_4, c32_0_4);
	full_adder ad32_0_5(a15_32, a16_32, a17_32, s32_0_5, c32_0_5);
	full_adder ad32_0_6(a18_32, a19_32, a20_32, s32_0_6, c32_0_6);
	full_adder ad32_0_7(a21_32, a22_32, a23_32, s32_0_7, c32_0_7);
	full_adder ad32_0_8(a24_32, a25_32, a26_32, s32_0_8, c32_0_8);
	full_adder ad32_0_9(a27_32, a28_32, a29_32, s32_0_9, c32_0_9);
	half_adder ha32_0_10(a30_32, a31_32, s32_0_10, c32_0_10);
	full_adder ad33_0_0(a2_33, a3_33, a4_33, s33_0_0, c33_0_0);
	full_adder ad33_0_1(a5_33, a6_33, a7_33, s33_0_1, c33_0_1);
	full_adder ad33_0_2(a8_33, a9_33, a10_33, s33_0_2, c33_0_2);
	full_adder ad33_0_3(a11_33, a12_33, a13_33, s33_0_3, c33_0_3);
	full_adder ad33_0_4(a14_33, a15_33, a16_33, s33_0_4, c33_0_4);
	full_adder ad33_0_5(a17_33, a18_33, a19_33, s33_0_5, c33_0_5);
	full_adder ad33_0_6(a20_33, a21_33, a22_33, s33_0_6, c33_0_6);
	full_adder ad33_0_7(a23_33, a24_33, a25_33, s33_0_7, c33_0_7);
	full_adder ad33_0_8(a26_33, a27_33, a28_33, s33_0_8, c33_0_8);
	full_adder ad33_0_9(a29_33, a30_33, a31_33, s33_0_9, c33_0_9);
	full_adder ad34_0_0(a3_34, a4_34, a5_34, s34_0_0, c34_0_0);
	full_adder ad34_0_1(a6_34, a7_34, a8_34, s34_0_1, c34_0_1);
	full_adder ad34_0_2(a9_34, a10_34, a11_34, s34_0_2, c34_0_2);
	full_adder ad34_0_3(a12_34, a13_34, a14_34, s34_0_3, c34_0_3);
	full_adder ad34_0_4(a15_34, a16_34, a17_34, s34_0_4, c34_0_4);
	full_adder ad34_0_5(a18_34, a19_34, a20_34, s34_0_5, c34_0_5);
	full_adder ad34_0_6(a21_34, a22_34, a23_34, s34_0_6, c34_0_6);
	full_adder ad34_0_7(a24_34, a25_34, a26_34, s34_0_7, c34_0_7);
	full_adder ad34_0_8(a27_34, a28_34, a29_34, s34_0_8, c34_0_8);
	half_adder ha34_0_9(a30_34, a31_34, s34_0_9, c34_0_9);
	full_adder ad35_0_0(a4_35, a5_35, a6_35, s35_0_0, c35_0_0);
	full_adder ad35_0_1(a7_35, a8_35, a9_35, s35_0_1, c35_0_1);
	full_adder ad35_0_2(a10_35, a11_35, a12_35, s35_0_2, c35_0_2);
	full_adder ad35_0_3(a13_35, a14_35, a15_35, s35_0_3, c35_0_3);
	full_adder ad35_0_4(a16_35, a17_35, a18_35, s35_0_4, c35_0_4);
	full_adder ad35_0_5(a19_35, a20_35, a21_35, s35_0_5, c35_0_5);
	full_adder ad35_0_6(a22_35, a23_35, a24_35, s35_0_6, c35_0_6);
	full_adder ad35_0_7(a25_35, a26_35, a27_35, s35_0_7, c35_0_7);
	full_adder ad35_0_8(a28_35, a29_35, a30_35, s35_0_8, c35_0_8);
	full_adder ad36_0_0(a5_36, a6_36, a7_36, s36_0_0, c36_0_0);
	full_adder ad36_0_1(a8_36, a9_36, a10_36, s36_0_1, c36_0_1);
	full_adder ad36_0_2(a11_36, a12_36, a13_36, s36_0_2, c36_0_2);
	full_adder ad36_0_3(a14_36, a15_36, a16_36, s36_0_3, c36_0_3);
	full_adder ad36_0_4(a17_36, a18_36, a19_36, s36_0_4, c36_0_4);
	full_adder ad36_0_5(a20_36, a21_36, a22_36, s36_0_5, c36_0_5);
	full_adder ad36_0_6(a23_36, a24_36, a25_36, s36_0_6, c36_0_6);
	full_adder ad36_0_7(a26_36, a27_36, a28_36, s36_0_7, c36_0_7);
	full_adder ad36_0_8(a29_36, a30_36, a31_36, s36_0_8, c36_0_8);
	full_adder ad37_0_0(a6_37, a7_37, a8_37, s37_0_0, c37_0_0);
	full_adder ad37_0_1(a9_37, a10_37, a11_37, s37_0_1, c37_0_1);
	full_adder ad37_0_2(a12_37, a13_37, a14_37, s37_0_2, c37_0_2);
	full_adder ad37_0_3(a15_37, a16_37, a17_37, s37_0_3, c37_0_3);
	full_adder ad37_0_4(a18_37, a19_37, a20_37, s37_0_4, c37_0_4);
	full_adder ad37_0_5(a21_37, a22_37, a23_37, s37_0_5, c37_0_5);
	full_adder ad37_0_6(a24_37, a25_37, a26_37, s37_0_6, c37_0_6);
	full_adder ad37_0_7(a27_37, a28_37, a29_37, s37_0_7, c37_0_7);
	half_adder ha37_0_8(a30_37, a31_37, s37_0_8, c37_0_8);
	full_adder ad38_0_0(a7_38, a8_38, a9_38, s38_0_0, c38_0_0);
	full_adder ad38_0_1(a10_38, a11_38, a12_38, s38_0_1, c38_0_1);
	full_adder ad38_0_2(a13_38, a14_38, a15_38, s38_0_2, c38_0_2);
	full_adder ad38_0_3(a16_38, a17_38, a18_38, s38_0_3, c38_0_3);
	full_adder ad38_0_4(a19_38, a20_38, a21_38, s38_0_4, c38_0_4);
	full_adder ad38_0_5(a22_38, a23_38, a24_38, s38_0_5, c38_0_5);
	full_adder ad38_0_6(a25_38, a26_38, a27_38, s38_0_6, c38_0_6);
	full_adder ad38_0_7(a28_38, a29_38, a30_38, s38_0_7, c38_0_7);
	full_adder ad39_0_0(a8_39, a9_39, a10_39, s39_0_0, c39_0_0);
	full_adder ad39_0_1(a11_39, a12_39, a13_39, s39_0_1, c39_0_1);
	full_adder ad39_0_2(a14_39, a15_39, a16_39, s39_0_2, c39_0_2);
	full_adder ad39_0_3(a17_39, a18_39, a19_39, s39_0_3, c39_0_3);
	full_adder ad39_0_4(a20_39, a21_39, a22_39, s39_0_4, c39_0_4);
	full_adder ad39_0_5(a23_39, a24_39, a25_39, s39_0_5, c39_0_5);
	full_adder ad39_0_6(a26_39, a27_39, a28_39, s39_0_6, c39_0_6);
	full_adder ad39_0_7(a29_39, a30_39, a31_39, s39_0_7, c39_0_7);
	full_adder ad40_0_0(a9_40, a10_40, a11_40, s40_0_0, c40_0_0);
	full_adder ad40_0_1(a12_40, a13_40, a14_40, s40_0_1, c40_0_1);
	full_adder ad40_0_2(a15_40, a16_40, a17_40, s40_0_2, c40_0_2);
	full_adder ad40_0_3(a18_40, a19_40, a20_40, s40_0_3, c40_0_3);
	full_adder ad40_0_4(a21_40, a22_40, a23_40, s40_0_4, c40_0_4);
	full_adder ad40_0_5(a24_40, a25_40, a26_40, s40_0_5, c40_0_5);
	full_adder ad40_0_6(a27_40, a28_40, a29_40, s40_0_6, c40_0_6);
	half_adder ha40_0_7(a30_40, a31_40, s40_0_7, c40_0_7);
	full_adder ad41_0_0(a10_41, a11_41, a12_41, s41_0_0, c41_0_0);
	full_adder ad41_0_1(a13_41, a14_41, a15_41, s41_0_1, c41_0_1);
	full_adder ad41_0_2(a16_41, a17_41, a18_41, s41_0_2, c41_0_2);
	full_adder ad41_0_3(a19_41, a20_41, a21_41, s41_0_3, c41_0_3);
	full_adder ad41_0_4(a22_41, a23_41, a24_41, s41_0_4, c41_0_4);
	full_adder ad41_0_5(a25_41, a26_41, a27_41, s41_0_5, c41_0_5);
	full_adder ad41_0_6(a28_41, a29_41, a30_41, s41_0_6, c41_0_6);
	full_adder ad42_0_0(a11_42, a12_42, a13_42, s42_0_0, c42_0_0);
	full_adder ad42_0_1(a14_42, a15_42, a16_42, s42_0_1, c42_0_1);
	full_adder ad42_0_2(a17_42, a18_42, a19_42, s42_0_2, c42_0_2);
	full_adder ad42_0_3(a20_42, a21_42, a22_42, s42_0_3, c42_0_3);
	full_adder ad42_0_4(a23_42, a24_42, a25_42, s42_0_4, c42_0_4);
	full_adder ad42_0_5(a26_42, a27_42, a28_42, s42_0_5, c42_0_5);
	full_adder ad42_0_6(a29_42, a30_42, a31_42, s42_0_6, c42_0_6);
	full_adder ad43_0_0(a12_43, a13_43, a14_43, s43_0_0, c43_0_0);
	full_adder ad43_0_1(a15_43, a16_43, a17_43, s43_0_1, c43_0_1);
	full_adder ad43_0_2(a18_43, a19_43, a20_43, s43_0_2, c43_0_2);
	full_adder ad43_0_3(a21_43, a22_43, a23_43, s43_0_3, c43_0_3);
	full_adder ad43_0_4(a24_43, a25_43, a26_43, s43_0_4, c43_0_4);
	full_adder ad43_0_5(a27_43, a28_43, a29_43, s43_0_5, c43_0_5);
	half_adder ha43_0_6(a30_43, a31_43, s43_0_6, c43_0_6);
	full_adder ad44_0_0(a13_44, a14_44, a15_44, s44_0_0, c44_0_0);
	full_adder ad44_0_1(a16_44, a17_44, a18_44, s44_0_1, c44_0_1);
	full_adder ad44_0_2(a19_44, a20_44, a21_44, s44_0_2, c44_0_2);
	full_adder ad44_0_3(a22_44, a23_44, a24_44, s44_0_3, c44_0_3);
	full_adder ad44_0_4(a25_44, a26_44, a27_44, s44_0_4, c44_0_4);
	full_adder ad44_0_5(a28_44, a29_44, a30_44, s44_0_5, c44_0_5);
	full_adder ad45_0_0(a14_45, a15_45, a16_45, s45_0_0, c45_0_0);
	full_adder ad45_0_1(a17_45, a18_45, a19_45, s45_0_1, c45_0_1);
	full_adder ad45_0_2(a20_45, a21_45, a22_45, s45_0_2, c45_0_2);
	full_adder ad45_0_3(a23_45, a24_45, a25_45, s45_0_3, c45_0_3);
	full_adder ad45_0_4(a26_45, a27_45, a28_45, s45_0_4, c45_0_4);
	full_adder ad45_0_5(a29_45, a30_45, a31_45, s45_0_5, c45_0_5);
	full_adder ad46_0_0(a15_46, a16_46, a17_46, s46_0_0, c46_0_0);
	full_adder ad46_0_1(a18_46, a19_46, a20_46, s46_0_1, c46_0_1);
	full_adder ad46_0_2(a21_46, a22_46, a23_46, s46_0_2, c46_0_2);
	full_adder ad46_0_3(a24_46, a25_46, a26_46, s46_0_3, c46_0_3);
	full_adder ad46_0_4(a27_46, a28_46, a29_46, s46_0_4, c46_0_4);
	half_adder ha46_0_5(a30_46, a31_46, s46_0_5, c46_0_5);
	full_adder ad47_0_0(a16_47, a17_47, a18_47, s47_0_0, c47_0_0);
	full_adder ad47_0_1(a19_47, a20_47, a21_47, s47_0_1, c47_0_1);
	full_adder ad47_0_2(a22_47, a23_47, a24_47, s47_0_2, c47_0_2);
	full_adder ad47_0_3(a25_47, a26_47, a27_47, s47_0_3, c47_0_3);
	full_adder ad47_0_4(a28_47, a29_47, a30_47, s47_0_4, c47_0_4);
	full_adder ad48_0_0(a17_48, a18_48, a19_48, s48_0_0, c48_0_0);
	full_adder ad48_0_1(a20_48, a21_48, a22_48, s48_0_1, c48_0_1);
	full_adder ad48_0_2(a23_48, a24_48, a25_48, s48_0_2, c48_0_2);
	full_adder ad48_0_3(a26_48, a27_48, a28_48, s48_0_3, c48_0_3);
	full_adder ad48_0_4(a29_48, a30_48, a31_48, s48_0_4, c48_0_4);
	full_adder ad49_0_0(a18_49, a19_49, a20_49, s49_0_0, c49_0_0);
	full_adder ad49_0_1(a21_49, a22_49, a23_49, s49_0_1, c49_0_1);
	full_adder ad49_0_2(a24_49, a25_49, a26_49, s49_0_2, c49_0_2);
	full_adder ad49_0_3(a27_49, a28_49, a29_49, s49_0_3, c49_0_3);
	half_adder ha49_0_4(a30_49, a31_49, s49_0_4, c49_0_4);
	full_adder ad50_0_0(a19_50, a20_50, a21_50, s50_0_0, c50_0_0);
	full_adder ad50_0_1(a22_50, a23_50, a24_50, s50_0_1, c50_0_1);
	full_adder ad50_0_2(a25_50, a26_50, a27_50, s50_0_2, c50_0_2);
	full_adder ad50_0_3(a28_50, a29_50, a30_50, s50_0_3, c50_0_3);
	full_adder ad51_0_0(a20_51, a21_51, a22_51, s51_0_0, c51_0_0);
	full_adder ad51_0_1(a23_51, a24_51, a25_51, s51_0_1, c51_0_1);
	full_adder ad51_0_2(a26_51, a27_51, a28_51, s51_0_2, c51_0_2);
	full_adder ad51_0_3(a29_51, a30_51, a31_51, s51_0_3, c51_0_3);
	full_adder ad52_0_0(a21_52, a22_52, a23_52, s52_0_0, c52_0_0);
	full_adder ad52_0_1(a24_52, a25_52, a26_52, s52_0_1, c52_0_1);
	full_adder ad52_0_2(a27_52, a28_52, a29_52, s52_0_2, c52_0_2);
	half_adder ha52_0_3(a30_52, a31_52, s52_0_3, c52_0_3);
	full_adder ad53_0_0(a22_53, a23_53, a24_53, s53_0_0, c53_0_0);
	full_adder ad53_0_1(a25_53, a26_53, a27_53, s53_0_1, c53_0_1);
	full_adder ad53_0_2(a28_53, a29_53, a30_53, s53_0_2, c53_0_2);
	full_adder ad54_0_0(a23_54, a24_54, a25_54, s54_0_0, c54_0_0);
	full_adder ad54_0_1(a26_54, a27_54, a28_54, s54_0_1, c54_0_1);
	full_adder ad54_0_2(a29_54, a30_54, a31_54, s54_0_2, c54_0_2);
	full_adder ad55_0_0(a24_55, a25_55, a26_55, s55_0_0, c55_0_0);
	full_adder ad55_0_1(a27_55, a28_55, a29_55, s55_0_1, c55_0_1);
	half_adder ha55_0_2(a30_55, a31_55, s55_0_2, c55_0_2);
	full_adder ad56_0_0(a25_56, a26_56, a27_56, s56_0_0, c56_0_0);
	full_adder ad56_0_1(a28_56, a29_56, a30_56, s56_0_1, c56_0_1);
	full_adder ad57_0_0(a26_57, a27_57, a28_57, s57_0_0, c57_0_0);
	full_adder ad57_0_1(a29_57, a30_57, a31_57, s57_0_1, c57_0_1);
	full_adder ad58_0_0(a27_58, a28_58, a29_58, s58_0_0, c58_0_0);
	half_adder ha58_0_1(a30_58, a31_58, s58_0_1, c58_0_1);
	full_adder ad59_0_0(a28_59, a29_59, a30_59, s59_0_0, c59_0_0);
	full_adder ad60_0_0(a29_60, a30_60, a31_60, s60_0_0, c60_0_0);
	half_adder ha61_0_0(a30_61, a31_61, s61_0_0, c61_0_0);

	half_adder ha2_1_0(c1_0_0, s2_0_0, s2_1_0, c2_1_0);
	full_adder ad3_1_0(c2_0_0, s3_0_0, a3_3, s3_1_0, c3_1_0);
	full_adder ad4_1_0(c3_0_0, s4_0_0, s4_0_1, s4_1_0, c4_1_0);
	full_adder ad5_1_0(c4_0_0, c4_0_1, s5_0_0, s5_1_0, c5_1_0);
	full_adder ad6_1_0(c5_0_0, c5_0_1, s6_0_0, s6_1_0, c6_1_0);
	half_adder ha6_1_1(s6_0_1, a6_6, s6_1_1, c6_1_1);
	full_adder ad7_1_0(c6_0_0, c6_0_1, s7_0_0, s7_1_0, c7_1_0);
	half_adder ha7_1_1(s7_0_1, s7_0_2, s7_1_1, c7_1_1);
	full_adder ad8_1_0(c7_0_0, c7_0_1, c7_0_2, s8_1_0, c8_1_0);
	full_adder ad8_1_1(s8_0_0, s8_0_1, s8_0_2, s8_1_1, c8_1_1);
	full_adder ad9_1_0(c8_0_0, c8_0_1, c8_0_2, s9_1_0, c9_1_0);
	full_adder ad9_1_1(s9_0_0, s9_0_1, s9_0_2, s9_1_1, c9_1_1);
	full_adder ad10_1_0(c9_0_0, c9_0_1, c9_0_2, s10_1_0, c10_1_0);
	full_adder ad10_1_1(s10_0_0, s10_0_1, s10_0_2, s10_1_1, c10_1_1);
	full_adder ad11_1_0(c10_0_0, c10_0_1, c10_0_2, s11_1_0, c11_1_0);
	full_adder ad11_1_1(c10_0_3, s11_0_0, s11_0_1, s11_1_1, c11_1_1);
	half_adder ha11_1_2(s11_0_2, s11_0_3, s11_1_2, c11_1_2);
	full_adder ad12_1_0(c11_0_0, c11_0_1, c11_0_2, s12_1_0, c12_1_0);
	full_adder ad12_1_1(c11_0_3, s12_0_0, s12_0_1, s12_1_1, c12_1_1);
	full_adder ad12_1_2(s12_0_2, s12_0_3, a12_12, s12_1_2, c12_1_2);
	full_adder ad13_1_0(c12_0_0, c12_0_1, c12_0_2, s13_1_0, c13_1_0);
	full_adder ad13_1_1(c12_0_3, s13_0_0, s13_0_1, s13_1_1, c13_1_1);
	full_adder ad13_1_2(s13_0_2, s13_0_3, s13_0_4, s13_1_2, c13_1_2);
	full_adder ad14_1_0(c13_0_0, c13_0_1, c13_0_2, s14_1_0, c14_1_0);
	full_adder ad14_1_1(c13_0_3, c13_0_4, s14_0_0, s14_1_1, c14_1_1);
	full_adder ad14_1_2(s14_0_1, s14_0_2, s14_0_3, s14_1_2, c14_1_2);
	full_adder ad15_1_0(c14_0_0, c14_0_1, c14_0_2, s15_1_0, c15_1_0);
	full_adder ad15_1_1(c14_0_3, c14_0_4, s15_0_0, s15_1_1, c15_1_1);
	full_adder ad15_1_2(s15_0_1, s15_0_2, s15_0_3, s15_1_2, c15_1_2);
	half_adder ha15_1_3(s15_0_4, a15_15, s15_1_3, c15_1_3);
	full_adder ad16_1_0(c15_0_0, c15_0_1, c15_0_2, s16_1_0, c16_1_0);
	full_adder ad16_1_1(c15_0_3, c15_0_4, s16_0_0, s16_1_1, c16_1_1);
	full_adder ad16_1_2(s16_0_1, s16_0_2, s16_0_3, s16_1_2, c16_1_2);
	half_adder ha16_1_3(s16_0_4, s16_0_5, s16_1_3, c16_1_3);
	full_adder ad17_1_0(c16_0_0, c16_0_1, c16_0_2, s17_1_0, c17_1_0);
	full_adder ad17_1_1(c16_0_3, c16_0_4, c16_0_5, s17_1_1, c17_1_1);
	full_adder ad17_1_2(s17_0_0, s17_0_1, s17_0_2, s17_1_2, c17_1_2);
	full_adder ad17_1_3(s17_0_3, s17_0_4, s17_0_5, s17_1_3, c17_1_3);
	full_adder ad18_1_0(c17_0_0, c17_0_1, c17_0_2, s18_1_0, c18_1_0);
	full_adder ad18_1_1(c17_0_3, c17_0_4, c17_0_5, s18_1_1, c18_1_1);
	full_adder ad18_1_2(s18_0_0, s18_0_1, s18_0_2, s18_1_2, c18_1_2);
	full_adder ad18_1_3(s18_0_3, s18_0_4, s18_0_5, s18_1_3, c18_1_3);
	full_adder ad19_1_0(c18_0_0, c18_0_1, c18_0_2, s19_1_0, c19_1_0);
	full_adder ad19_1_1(c18_0_3, c18_0_4, c18_0_5, s19_1_1, c19_1_1);
	full_adder ad19_1_2(s19_0_0, s19_0_1, s19_0_2, s19_1_2, c19_1_2);
	full_adder ad19_1_3(s19_0_3, s19_0_4, s19_0_5, s19_1_3, c19_1_3);
	full_adder ad20_1_0(c19_0_0, c19_0_1, c19_0_2, s20_1_0, c20_1_0);
	full_adder ad20_1_1(c19_0_3, c19_0_4, c19_0_5, s20_1_1, c20_1_1);
	full_adder ad20_1_2(c19_0_6, s20_0_0, s20_0_1, s20_1_2, c20_1_2);
	full_adder ad20_1_3(s20_0_2, s20_0_3, s20_0_4, s20_1_3, c20_1_3);
	half_adder ha20_1_4(s20_0_5, s20_0_6, s20_1_4, c20_1_4);
	full_adder ad21_1_0(c20_0_0, c20_0_1, c20_0_2, s21_1_0, c21_1_0);
	full_adder ad21_1_1(c20_0_3, c20_0_4, c20_0_5, s21_1_1, c21_1_1);
	full_adder ad21_1_2(c20_0_6, s21_0_0, s21_0_1, s21_1_2, c21_1_2);
	full_adder ad21_1_3(s21_0_2, s21_0_3, s21_0_4, s21_1_3, c21_1_3);
	full_adder ad21_1_4(s21_0_5, s21_0_6, a21_21, s21_1_4, c21_1_4);
	full_adder ad22_1_0(c21_0_0, c21_0_1, c21_0_2, s22_1_0, c22_1_0);
	full_adder ad22_1_1(c21_0_3, c21_0_4, c21_0_5, s22_1_1, c22_1_1);
	full_adder ad22_1_2(c21_0_6, s22_0_0, s22_0_1, s22_1_2, c22_1_2);
	full_adder ad22_1_3(s22_0_2, s22_0_3, s22_0_4, s22_1_3, c22_1_3);
	full_adder ad22_1_4(s22_0_5, s22_0_6, s22_0_7, s22_1_4, c22_1_4);
	full_adder ad23_1_0(c22_0_0, c22_0_1, c22_0_2, s23_1_0, c23_1_0);
	full_adder ad23_1_1(c22_0_3, c22_0_4, c22_0_5, s23_1_1, c23_1_1);
	full_adder ad23_1_2(c22_0_6, c22_0_7, s23_0_0, s23_1_2, c23_1_2);
	full_adder ad23_1_3(s23_0_1, s23_0_2, s23_0_3, s23_1_3, c23_1_3);
	full_adder ad23_1_4(s23_0_4, s23_0_5, s23_0_6, s23_1_4, c23_1_4);
	full_adder ad24_1_0(c23_0_0, c23_0_1, c23_0_2, s24_1_0, c24_1_0);
	full_adder ad24_1_1(c23_0_3, c23_0_4, c23_0_5, s24_1_1, c24_1_1);
	full_adder ad24_1_2(c23_0_6, c23_0_7, s24_0_0, s24_1_2, c24_1_2);
	full_adder ad24_1_3(s24_0_1, s24_0_2, s24_0_3, s24_1_3, c24_1_3);
	full_adder ad24_1_4(s24_0_4, s24_0_5, s24_0_6, s24_1_4, c24_1_4);
	half_adder ha24_1_5(s24_0_7, a24_24, s24_1_5, c24_1_5);
	full_adder ad25_1_0(c24_0_0, c24_0_1, c24_0_2, s25_1_0, c25_1_0);
	full_adder ad25_1_1(c24_0_3, c24_0_4, c24_0_5, s25_1_1, c25_1_1);
	full_adder ad25_1_2(c24_0_6, c24_0_7, s25_0_0, s25_1_2, c25_1_2);
	full_adder ad25_1_3(s25_0_1, s25_0_2, s25_0_3, s25_1_3, c25_1_3);
	full_adder ad25_1_4(s25_0_4, s25_0_5, s25_0_6, s25_1_4, c25_1_4);
	half_adder ha25_1_5(s25_0_7, s25_0_8, s25_1_5, c25_1_5);
	full_adder ad26_1_0(c25_0_0, c25_0_1, c25_0_2, s26_1_0, c26_1_0);
	full_adder ad26_1_1(c25_0_3, c25_0_4, c25_0_5, s26_1_1, c26_1_1);
	full_adder ad26_1_2(c25_0_6, c25_0_7, c25_0_8, s26_1_2, c26_1_2);
	full_adder ad26_1_3(s26_0_0, s26_0_1, s26_0_2, s26_1_3, c26_1_3);
	full_adder ad26_1_4(s26_0_3, s26_0_4, s26_0_5, s26_1_4, c26_1_4);
	full_adder ad26_1_5(s26_0_6, s26_0_7, s26_0_8, s26_1_5, c26_1_5);
	full_adder ad27_1_0(c26_0_0, c26_0_1, c26_0_2, s27_1_0, c27_1_0);
	full_adder ad27_1_1(c26_0_3, c26_0_4, c26_0_5, s27_1_1, c27_1_1);
	full_adder ad27_1_2(c26_0_6, c26_0_7, c26_0_8, s27_1_2, c27_1_2);
	full_adder ad27_1_3(s27_0_0, s27_0_1, s27_0_2, s27_1_3, c27_1_3);
	full_adder ad27_1_4(s27_0_3, s27_0_4, s27_0_5, s27_1_4, c27_1_4);
	full_adder ad27_1_5(s27_0_6, s27_0_7, s27_0_8, s27_1_5, c27_1_5);
	full_adder ad28_1_0(c27_0_0, c27_0_1, c27_0_2, s28_1_0, c28_1_0);
	full_adder ad28_1_1(c27_0_3, c27_0_4, c27_0_5, s28_1_1, c28_1_1);
	full_adder ad28_1_2(c27_0_6, c27_0_7, c27_0_8, s28_1_2, c28_1_2);
	full_adder ad28_1_3(s28_0_0, s28_0_1, s28_0_2, s28_1_3, c28_1_3);
	full_adder ad28_1_4(s28_0_3, s28_0_4, s28_0_5, s28_1_4, c28_1_4);
	full_adder ad28_1_5(s28_0_6, s28_0_7, s28_0_8, s28_1_5, c28_1_5);
	full_adder ad29_1_0(c28_0_0, c28_0_1, c28_0_2, s29_1_0, c29_1_0);
	full_adder ad29_1_1(c28_0_3, c28_0_4, c28_0_5, s29_1_1, c29_1_1);
	full_adder ad29_1_2(c28_0_6, c28_0_7, c28_0_8, s29_1_2, c29_1_2);
	full_adder ad29_1_3(c28_0_9, s29_0_0, s29_0_1, s29_1_3, c29_1_3);
	full_adder ad29_1_4(s29_0_2, s29_0_3, s29_0_4, s29_1_4, c29_1_4);
	full_adder ad29_1_5(s29_0_5, s29_0_6, s29_0_7, s29_1_5, c29_1_5);
	half_adder ha29_1_6(s29_0_8, s29_0_9, s29_1_6, c29_1_6);
	full_adder ad30_1_0(c29_0_0, c29_0_1, c29_0_2, s30_1_0, c30_1_0);
	full_adder ad30_1_1(c29_0_3, c29_0_4, c29_0_5, s30_1_1, c30_1_1);
	full_adder ad30_1_2(c29_0_6, c29_0_7, c29_0_8, s30_1_2, c30_1_2);
	full_adder ad30_1_3(c29_0_9, s30_0_0, s30_0_1, s30_1_3, c30_1_3);
	full_adder ad30_1_4(s30_0_2, s30_0_3, s30_0_4, s30_1_4, c30_1_4);
	full_adder ad30_1_5(s30_0_5, s30_0_6, s30_0_7, s30_1_5, c30_1_5);
	full_adder ad30_1_6(s30_0_8, s30_0_9, a30_30, s30_1_6, c30_1_6);
	full_adder ad31_1_0(c30_0_0, c30_0_1, c30_0_2, s31_1_0, c31_1_0);
	full_adder ad31_1_1(c30_0_3, c30_0_4, c30_0_5, s31_1_1, c31_1_1);
	full_adder ad31_1_2(c30_0_6, c30_0_7, c30_0_8, s31_1_2, c31_1_2);
	full_adder ad31_1_3(c30_0_9, s31_0_0, s31_0_1, s31_1_3, c31_1_3);
	full_adder ad31_1_4(s31_0_2, s31_0_3, s31_0_4, s31_1_4, c31_1_4);
	full_adder ad31_1_5(s31_0_5, s31_0_6, s31_0_7, s31_1_5, c31_1_5);
	full_adder ad31_1_6(s31_0_8, s31_0_9, s31_0_10, s31_1_6, c31_1_6);
	full_adder ad32_1_0(c31_0_0, c31_0_1, c31_0_2, s32_1_0, c32_1_0);
	full_adder ad32_1_1(c31_0_3, c31_0_4, c31_0_5, s32_1_1, c32_1_1);
	full_adder ad32_1_2(c31_0_6, c31_0_7, c31_0_8, s32_1_2, c32_1_2);
	full_adder ad32_1_3(c31_0_9, c31_0_10, s32_0_0, s32_1_3, c32_1_3);
	full_adder ad32_1_4(s32_0_1, s32_0_2, s32_0_3, s32_1_4, c32_1_4);
	full_adder ad32_1_5(s32_0_4, s32_0_5, s32_0_6, s32_1_5, c32_1_5);
	full_adder ad32_1_6(s32_0_7, s32_0_8, s32_0_9, s32_1_6, c32_1_6);
	full_adder ad33_1_0(c32_0_0, c32_0_1, c32_0_2, s33_1_0, c33_1_0);
	full_adder ad33_1_1(c32_0_3, c32_0_4, c32_0_5, s33_1_1, c33_1_1);
	full_adder ad33_1_2(c32_0_6, c32_0_7, c32_0_8, s33_1_2, c33_1_2);
	full_adder ad33_1_3(c32_0_9, c32_0_10, s33_0_0, s33_1_3, c33_1_3);
	full_adder ad33_1_4(s33_0_1, s33_0_2, s33_0_3, s33_1_4, c33_1_4);
	full_adder ad33_1_5(s33_0_4, s33_0_5, s33_0_6, s33_1_5, c33_1_5);
	full_adder ad33_1_6(s33_0_7, s33_0_8, s33_0_9, s33_1_6, c33_1_6);
	full_adder ad34_1_0(c33_0_0, c33_0_1, c33_0_2, s34_1_0, c34_1_0);
	full_adder ad34_1_1(c33_0_3, c33_0_4, c33_0_5, s34_1_1, c34_1_1);
	full_adder ad34_1_2(c33_0_6, c33_0_7, c33_0_8, s34_1_2, c34_1_2);
	full_adder ad34_1_3(c33_0_9, s34_0_0, s34_0_1, s34_1_3, c34_1_3);
	full_adder ad34_1_4(s34_0_2, s34_0_3, s34_0_4, s34_1_4, c34_1_4);
	full_adder ad34_1_5(s34_0_5, s34_0_6, s34_0_7, s34_1_5, c34_1_5);
	half_adder ha34_1_6(s34_0_8, s34_0_9, s34_1_6, c34_1_6);
	full_adder ad35_1_0(c34_0_0, c34_0_1, c34_0_2, s35_1_0, c35_1_0);
	full_adder ad35_1_1(c34_0_3, c34_0_4, c34_0_5, s35_1_1, c35_1_1);
	full_adder ad35_1_2(c34_0_6, c34_0_7, c34_0_8, s35_1_2, c35_1_2);
	full_adder ad35_1_3(c34_0_9, s35_0_0, s35_0_1, s35_1_3, c35_1_3);
	full_adder ad35_1_4(s35_0_2, s35_0_3, s35_0_4, s35_1_4, c35_1_4);
	full_adder ad35_1_5(s35_0_5, s35_0_6, s35_0_7, s35_1_5, c35_1_5);
	half_adder ha35_1_6(s35_0_8, a31_35, s35_1_6, c35_1_6);
	full_adder ad36_1_0(c35_0_0, c35_0_1, c35_0_2, s36_1_0, c36_1_0);
	full_adder ad36_1_1(c35_0_3, c35_0_4, c35_0_5, s36_1_1, c36_1_1);
	full_adder ad36_1_2(c35_0_6, c35_0_7, c35_0_8, s36_1_2, c36_1_2);
	full_adder ad36_1_3(s36_0_0, s36_0_1, s36_0_2, s36_1_3, c36_1_3);
	full_adder ad36_1_4(s36_0_3, s36_0_4, s36_0_5, s36_1_4, c36_1_4);
	full_adder ad36_1_5(s36_0_6, s36_0_7, s36_0_8, s36_1_5, c36_1_5);
	full_adder ad37_1_0(c36_0_0, c36_0_1, c36_0_2, s37_1_0, c37_1_0);
	full_adder ad37_1_1(c36_0_3, c36_0_4, c36_0_5, s37_1_1, c37_1_1);
	full_adder ad37_1_2(c36_0_6, c36_0_7, c36_0_8, s37_1_2, c37_1_2);
	full_adder ad37_1_3(s37_0_0, s37_0_1, s37_0_2, s37_1_3, c37_1_3);
	full_adder ad37_1_4(s37_0_3, s37_0_4, s37_0_5, s37_1_4, c37_1_4);
	full_adder ad37_1_5(s37_0_6, s37_0_7, s37_0_8, s37_1_5, c37_1_5);
	full_adder ad38_1_0(c37_0_0, c37_0_1, c37_0_2, s38_1_0, c38_1_0);
	full_adder ad38_1_1(c37_0_3, c37_0_4, c37_0_5, s38_1_1, c38_1_1);
	full_adder ad38_1_2(c37_0_6, c37_0_7, c37_0_8, s38_1_2, c38_1_2);
	full_adder ad38_1_3(s38_0_0, s38_0_1, s38_0_2, s38_1_3, c38_1_3);
	full_adder ad38_1_4(s38_0_3, s38_0_4, s38_0_5, s38_1_4, c38_1_4);
	full_adder ad38_1_5(s38_0_6, s38_0_7, a31_38, s38_1_5, c38_1_5);
	full_adder ad39_1_0(c38_0_0, c38_0_1, c38_0_2, s39_1_0, c39_1_0);
	full_adder ad39_1_1(c38_0_3, c38_0_4, c38_0_5, s39_1_1, c39_1_1);
	full_adder ad39_1_2(c38_0_6, c38_0_7, s39_0_0, s39_1_2, c39_1_2);
	full_adder ad39_1_3(s39_0_1, s39_0_2, s39_0_3, s39_1_3, c39_1_3);
	full_adder ad39_1_4(s39_0_4, s39_0_5, s39_0_6, s39_1_4, c39_1_4);
	full_adder ad40_1_0(c39_0_0, c39_0_1, c39_0_2, s40_1_0, c40_1_0);
	full_adder ad40_1_1(c39_0_3, c39_0_4, c39_0_5, s40_1_1, c40_1_1);
	full_adder ad40_1_2(c39_0_6, c39_0_7, s40_0_0, s40_1_2, c40_1_2);
	full_adder ad40_1_3(s40_0_1, s40_0_2, s40_0_3, s40_1_3, c40_1_3);
	full_adder ad40_1_4(s40_0_4, s40_0_5, s40_0_6, s40_1_4, c40_1_4);
	full_adder ad41_1_0(c40_0_0, c40_0_1, c40_0_2, s41_1_0, c41_1_0);
	full_adder ad41_1_1(c40_0_3, c40_0_4, c40_0_5, s41_1_1, c41_1_1);
	full_adder ad41_1_2(c40_0_6, c40_0_7, s41_0_0, s41_1_2, c41_1_2);
	full_adder ad41_1_3(s41_0_1, s41_0_2, s41_0_3, s41_1_3, c41_1_3);
	full_adder ad41_1_4(s41_0_4, s41_0_5, s41_0_6, s41_1_4, c41_1_4);
	full_adder ad42_1_0(c41_0_0, c41_0_1, c41_0_2, s42_1_0, c42_1_0);
	full_adder ad42_1_1(c41_0_3, c41_0_4, c41_0_5, s42_1_1, c42_1_1);
	full_adder ad42_1_2(c41_0_6, s42_0_0, s42_0_1, s42_1_2, c42_1_2);
	full_adder ad42_1_3(s42_0_2, s42_0_3, s42_0_4, s42_1_3, c42_1_3);
	half_adder ha42_1_4(s42_0_5, s42_0_6, s42_1_4, c42_1_4);
	full_adder ad43_1_0(c42_0_0, c42_0_1, c42_0_2, s43_1_0, c43_1_0);
	full_adder ad43_1_1(c42_0_3, c42_0_4, c42_0_5, s43_1_1, c43_1_1);
	full_adder ad43_1_2(c42_0_6, s43_0_0, s43_0_1, s43_1_2, c43_1_2);
	full_adder ad43_1_3(s43_0_2, s43_0_3, s43_0_4, s43_1_3, c43_1_3);
	half_adder ha43_1_4(s43_0_5, s43_0_6, s43_1_4, c43_1_4);
	full_adder ad44_1_0(c43_0_0, c43_0_1, c43_0_2, s44_1_0, c44_1_0);
	full_adder ad44_1_1(c43_0_3, c43_0_4, c43_0_5, s44_1_1, c44_1_1);
	full_adder ad44_1_2(c43_0_6, s44_0_0, s44_0_1, s44_1_2, c44_1_2);
	full_adder ad44_1_3(s44_0_2, s44_0_3, s44_0_4, s44_1_3, c44_1_3);
	half_adder ha44_1_4(s44_0_5, a31_44, s44_1_4, c44_1_4);
	full_adder ad45_1_0(c44_0_0, c44_0_1, c44_0_2, s45_1_0, c45_1_0);
	full_adder ad45_1_1(c44_0_3, c44_0_4, c44_0_5, s45_1_1, c45_1_1);
	full_adder ad45_1_2(s45_0_0, s45_0_1, s45_0_2, s45_1_2, c45_1_2);
	full_adder ad45_1_3(s45_0_3, s45_0_4, s45_0_5, s45_1_3, c45_1_3);
	full_adder ad46_1_0(c45_0_0, c45_0_1, c45_0_2, s46_1_0, c46_1_0);
	full_adder ad46_1_1(c45_0_3, c45_0_4, c45_0_5, s46_1_1, c46_1_1);
	full_adder ad46_1_2(s46_0_0, s46_0_1, s46_0_2, s46_1_2, c46_1_2);
	full_adder ad46_1_3(s46_0_3, s46_0_4, s46_0_5, s46_1_3, c46_1_3);
	full_adder ad47_1_0(c46_0_0, c46_0_1, c46_0_2, s47_1_0, c47_1_0);
	full_adder ad47_1_1(c46_0_3, c46_0_4, c46_0_5, s47_1_1, c47_1_1);
	full_adder ad47_1_2(s47_0_0, s47_0_1, s47_0_2, s47_1_2, c47_1_2);
	full_adder ad47_1_3(s47_0_3, s47_0_4, a31_47, s47_1_3, c47_1_3);
	full_adder ad48_1_0(c47_0_0, c47_0_1, c47_0_2, s48_1_0, c48_1_0);
	full_adder ad48_1_1(c47_0_3, c47_0_4, s48_0_0, s48_1_1, c48_1_1);
	full_adder ad48_1_2(s48_0_1, s48_0_2, s48_0_3, s48_1_2, c48_1_2);
	full_adder ad49_1_0(c48_0_0, c48_0_1, c48_0_2, s49_1_0, c49_1_0);
	full_adder ad49_1_1(c48_0_3, c48_0_4, s49_0_0, s49_1_1, c49_1_1);
	full_adder ad49_1_2(s49_0_1, s49_0_2, s49_0_3, s49_1_2, c49_1_2);
	full_adder ad50_1_0(c49_0_0, c49_0_1, c49_0_2, s50_1_0, c50_1_0);
	full_adder ad50_1_1(c49_0_3, c49_0_4, s50_0_0, s50_1_1, c50_1_1);
	full_adder ad50_1_2(s50_0_1, s50_0_2, s50_0_3, s50_1_2, c50_1_2);
	full_adder ad51_1_0(c50_0_0, c50_0_1, c50_0_2, s51_1_0, c51_1_0);
	full_adder ad51_1_1(c50_0_3, s51_0_0, s51_0_1, s51_1_1, c51_1_1);
	half_adder ha51_1_2(s51_0_2, s51_0_3, s51_1_2, c51_1_2);
	full_adder ad52_1_0(c51_0_0, c51_0_1, c51_0_2, s52_1_0, c52_1_0);
	full_adder ad52_1_1(c51_0_3, s52_0_0, s52_0_1, s52_1_1, c52_1_1);
	half_adder ha52_1_2(s52_0_2, s52_0_3, s52_1_2, c52_1_2);
	full_adder ad53_1_0(c52_0_0, c52_0_1, c52_0_2, s53_1_0, c53_1_0);
	full_adder ad53_1_1(c52_0_3, s53_0_0, s53_0_1, s53_1_1, c53_1_1);
	half_adder ha53_1_2(s53_0_2, a31_53, s53_1_2, c53_1_2);
	full_adder ad54_1_0(c53_0_0, c53_0_1, c53_0_2, s54_1_0, c54_1_0);
	full_adder ad54_1_1(s54_0_0, s54_0_1, s54_0_2, s54_1_1, c54_1_1);
	full_adder ad55_1_0(c54_0_0, c54_0_1, c54_0_2, s55_1_0, c55_1_0);
	full_adder ad55_1_1(s55_0_0, s55_0_1, s55_0_2, s55_1_1, c55_1_1);
	full_adder ad56_1_0(c55_0_0, c55_0_1, c55_0_2, s56_1_0, c56_1_0);
	full_adder ad56_1_1(s56_0_0, s56_0_1, a31_56, s56_1_1, c56_1_1);
	full_adder ad57_1_0(c56_0_0, c56_0_1, s57_0_0, s57_1_0, c57_1_0);
	full_adder ad58_1_0(c57_0_0, c57_0_1, s58_0_0, s58_1_0, c58_1_0);
	full_adder ad59_1_0(c58_0_0, c58_0_1, s59_0_0, s59_1_0, c59_1_0);
	half_adder ha60_1_0(c59_0_0, s60_0_0, s60_1_0, c60_1_0);
	half_adder ha61_1_0(c60_0_0, s61_0_0, s61_1_0, c61_1_0);
	half_adder ha62_1_0(c61_0_0, a31_62, s62_1_0, c62_1_0);

	half_adder ha3_2_0(c2_1_0, s3_1_0, s3_2_0, c3_2_0);
	half_adder ha4_2_0(c3_1_0, s4_1_0, s4_2_0, c4_2_0);
	full_adder ad5_2_0(c4_1_0, s5_1_0, s5_0_1, s5_2_0, c5_2_0);
	full_adder ad6_2_0(c5_1_0, s6_1_0, s6_1_1, s6_2_0, c6_2_0);
	full_adder ad7_2_0(c6_1_0, c6_1_1, s7_1_0, s7_2_0, c7_2_0);
	full_adder ad8_2_0(c7_1_0, c7_1_1, s8_1_0, s8_2_0, c8_2_0);
	full_adder ad9_2_0(c8_1_0, c8_1_1, s9_1_0, s9_2_0, c9_2_0);
	half_adder ha9_2_1(s9_1_1, a9_9, s9_2_1, c9_2_1);
	full_adder ad10_2_0(c9_1_0, c9_1_1, s10_1_0, s10_2_0, c10_2_0);
	half_adder ha10_2_1(s10_1_1, s10_0_3, s10_2_1, c10_2_1);
	full_adder ad11_2_0(c10_1_0, c10_1_1, s11_1_0, s11_2_0, c11_2_0);
	half_adder ha11_2_1(s11_1_1, s11_1_2, s11_2_1, c11_2_1);
	full_adder ad12_2_0(c11_1_0, c11_1_1, c11_1_2, s12_2_0, c12_2_0);
	full_adder ad12_2_1(s12_1_0, s12_1_1, s12_1_2, s12_2_1, c12_2_1);
	full_adder ad13_2_0(c12_1_0, c12_1_1, c12_1_2, s13_2_0, c13_2_0);
	full_adder ad13_2_1(s13_1_0, s13_1_1, s13_1_2, s13_2_1, c13_2_1);
	full_adder ad14_2_0(c13_1_0, c13_1_1, c13_1_2, s14_2_0, c14_2_0);
	full_adder ad14_2_1(s14_1_0, s14_1_1, s14_1_2, s14_2_1, c14_2_1);
	full_adder ad15_2_0(c14_1_0, c14_1_1, c14_1_2, s15_2_0, c15_2_0);
	full_adder ad15_2_1(s15_1_0, s15_1_1, s15_1_2, s15_2_1, c15_2_1);
	full_adder ad16_2_0(c15_1_0, c15_1_1, c15_1_2, s16_2_0, c16_2_0);
	full_adder ad16_2_1(c15_1_3, s16_1_0, s16_1_1, s16_2_1, c16_2_1);
	half_adder ha16_2_2(s16_1_2, s16_1_3, s16_2_2, c16_2_2);
	full_adder ad17_2_0(c16_1_0, c16_1_1, c16_1_2, s17_2_0, c17_2_0);
	full_adder ad17_2_1(c16_1_3, s17_1_0, s17_1_1, s17_2_1, c17_2_1);
	half_adder ha17_2_2(s17_1_2, s17_1_3, s17_2_2, c17_2_2);
	full_adder ad18_2_0(c17_1_0, c17_1_1, c17_1_2, s18_2_0, c18_2_0);
	full_adder ad18_2_1(c17_1_3, s18_1_0, s18_1_1, s18_2_1, c18_2_1);
	full_adder ad18_2_2(s18_1_2, s18_1_3, a18_18, s18_2_2, c18_2_2);
	full_adder ad19_2_0(c18_1_0, c18_1_1, c18_1_2, s19_2_0, c19_2_0);
	full_adder ad19_2_1(c18_1_3, s19_1_0, s19_1_1, s19_2_1, c19_2_1);
	full_adder ad19_2_2(s19_1_2, s19_1_3, s19_0_6, s19_2_2, c19_2_2);
	full_adder ad20_2_0(c19_1_0, c19_1_1, c19_1_2, s20_2_0, c20_2_0);
	full_adder ad20_2_1(c19_1_3, s20_1_0, s20_1_1, s20_2_1, c20_2_1);
	full_adder ad20_2_2(s20_1_2, s20_1_3, s20_1_4, s20_2_2, c20_2_2);
	full_adder ad21_2_0(c20_1_0, c20_1_1, c20_1_2, s21_2_0, c21_2_0);
	full_adder ad21_2_1(c20_1_3, c20_1_4, s21_1_0, s21_2_1, c21_2_1);
	full_adder ad21_2_2(s21_1_1, s21_1_2, s21_1_3, s21_2_2, c21_2_2);
	full_adder ad22_2_0(c21_1_0, c21_1_1, c21_1_2, s22_2_0, c22_2_0);
	full_adder ad22_2_1(c21_1_3, c21_1_4, s22_1_0, s22_2_1, c22_2_1);
	full_adder ad22_2_2(s22_1_1, s22_1_2, s22_1_3, s22_2_2, c22_2_2);
	full_adder ad23_2_0(c22_1_0, c22_1_1, c22_1_2, s23_2_0, c23_2_0);
	full_adder ad23_2_1(c22_1_3, c22_1_4, s23_1_0, s23_2_1, c23_2_1);
	full_adder ad23_2_2(s23_1_1, s23_1_2, s23_1_3, s23_2_2, c23_2_2);
	half_adder ha23_2_3(s23_1_4, s23_0_7, s23_2_3, c23_2_3);
	full_adder ad24_2_0(c23_1_0, c23_1_1, c23_1_2, s24_2_0, c24_2_0);
	full_adder ad24_2_1(c23_1_3, c23_1_4, s24_1_0, s24_2_1, c24_2_1);
	full_adder ad24_2_2(s24_1_1, s24_1_2, s24_1_3, s24_2_2, c24_2_2);
	half_adder ha24_2_3(s24_1_4, s24_1_5, s24_2_3, c24_2_3);
	full_adder ad25_2_0(c24_1_0, c24_1_1, c24_1_2, s25_2_0, c25_2_0);
	full_adder ad25_2_1(c24_1_3, c24_1_4, c24_1_5, s25_2_1, c25_2_1);
	full_adder ad25_2_2(s25_1_0, s25_1_1, s25_1_2, s25_2_2, c25_2_2);
	full_adder ad25_2_3(s25_1_3, s25_1_4, s25_1_5, s25_2_3, c25_2_3);
	full_adder ad26_2_0(c25_1_0, c25_1_1, c25_1_2, s26_2_0, c26_2_0);
	full_adder ad26_2_1(c25_1_3, c25_1_4, c25_1_5, s26_2_1, c26_2_1);
	full_adder ad26_2_2(s26_1_0, s26_1_1, s26_1_2, s26_2_2, c26_2_2);
	full_adder ad26_2_3(s26_1_3, s26_1_4, s26_1_5, s26_2_3, c26_2_3);
	full_adder ad27_2_0(c26_1_0, c26_1_1, c26_1_2, s27_2_0, c27_2_0);
	full_adder ad27_2_1(c26_1_3, c26_1_4, c26_1_5, s27_2_1, c27_2_1);
	full_adder ad27_2_2(s27_1_0, s27_1_1, s27_1_2, s27_2_2, c27_2_2);
	full_adder ad27_2_3(s27_1_3, s27_1_4, s27_1_5, s27_2_3, c27_2_3);
	full_adder ad28_2_0(c27_1_0, c27_1_1, c27_1_2, s28_2_0, c28_2_0);
	full_adder ad28_2_1(c27_1_3, c27_1_4, c27_1_5, s28_2_1, c28_2_1);
	full_adder ad28_2_2(s28_1_0, s28_1_1, s28_1_2, s28_2_2, c28_2_2);
	full_adder ad28_2_3(s28_1_3, s28_1_4, s28_1_5, s28_2_3, c28_2_3);
	full_adder ad29_2_0(c28_1_0, c28_1_1, c28_1_2, s29_2_0, c29_2_0);
	full_adder ad29_2_1(c28_1_3, c28_1_4, c28_1_5, s29_2_1, c29_2_1);
	full_adder ad29_2_2(s29_1_0, s29_1_1, s29_1_2, s29_2_2, c29_2_2);
	full_adder ad29_2_3(s29_1_3, s29_1_4, s29_1_5, s29_2_3, c29_2_3);
	full_adder ad30_2_0(c29_1_0, c29_1_1, c29_1_2, s30_2_0, c30_2_0);
	full_adder ad30_2_1(c29_1_3, c29_1_4, c29_1_5, s30_2_1, c30_2_1);
	full_adder ad30_2_2(c29_1_6, s30_1_0, s30_1_1, s30_2_2, c30_2_2);
	full_adder ad30_2_3(s30_1_2, s30_1_3, s30_1_4, s30_2_3, c30_2_3);
	half_adder ha30_2_4(s30_1_5, s30_1_6, s30_2_4, c30_2_4);
	full_adder ad31_2_0(c30_1_0, c30_1_1, c30_1_2, s31_2_0, c31_2_0);
	full_adder ad31_2_1(c30_1_3, c30_1_4, c30_1_5, s31_2_1, c31_2_1);
	full_adder ad31_2_2(c30_1_6, s31_1_0, s31_1_1, s31_2_2, c31_2_2);
	full_adder ad31_2_3(s31_1_2, s31_1_3, s31_1_4, s31_2_3, c31_2_3);
	half_adder ha31_2_4(s31_1_5, s31_1_6, s31_2_4, c31_2_4);
	full_adder ad32_2_0(c31_1_0, c31_1_1, c31_1_2, s32_2_0, c32_2_0);
	full_adder ad32_2_1(c31_1_3, c31_1_4, c31_1_5, s32_2_1, c32_2_1);
	full_adder ad32_2_2(c31_1_6, s32_1_0, s32_1_1, s32_2_2, c32_2_2);
	full_adder ad32_2_3(s32_1_2, s32_1_3, s32_1_4, s32_2_3, c32_2_3);
	full_adder ad32_2_4(s32_1_5, s32_1_6, s32_0_10, s32_2_4, c32_2_4);
	full_adder ad33_2_0(c32_1_0, c32_1_1, c32_1_2, s33_2_0, c33_2_0);
	full_adder ad33_2_1(c32_1_3, c32_1_4, c32_1_5, s33_2_1, c33_2_1);
	full_adder ad33_2_2(c32_1_6, s33_1_0, s33_1_1, s33_2_2, c33_2_2);
	full_adder ad33_2_3(s33_1_2, s33_1_3, s33_1_4, s33_2_3, c33_2_3);
	half_adder ha33_2_4(s33_1_5, s33_1_6, s33_2_4, c33_2_4);
	full_adder ad34_2_0(c33_1_0, c33_1_1, c33_1_2, s34_2_0, c34_2_0);
	full_adder ad34_2_1(c33_1_3, c33_1_4, c33_1_5, s34_2_1, c34_2_1);
	full_adder ad34_2_2(c33_1_6, s34_1_0, s34_1_1, s34_2_2, c34_2_2);
	full_adder ad34_2_3(s34_1_2, s34_1_3, s34_1_4, s34_2_3, c34_2_3);
	half_adder ha34_2_4(s34_1_5, s34_1_6, s34_2_4, c34_2_4);
	full_adder ad35_2_0(c34_1_0, c34_1_1, c34_1_2, s35_2_0, c35_2_0);
	full_adder ad35_2_1(c34_1_3, c34_1_4, c34_1_5, s35_2_1, c35_2_1);
	full_adder ad35_2_2(c34_1_6, s35_1_0, s35_1_1, s35_2_2, c35_2_2);
	full_adder ad35_2_3(s35_1_2, s35_1_3, s35_1_4, s35_2_3, c35_2_3);
	half_adder ha35_2_4(s35_1_5, s35_1_6, s35_2_4, c35_2_4);
	full_adder ad36_2_0(c35_1_0, c35_1_1, c35_1_2, s36_2_0, c36_2_0);
	full_adder ad36_2_1(c35_1_3, c35_1_4, c35_1_5, s36_2_1, c36_2_1);
	full_adder ad36_2_2(c35_1_6, s36_1_0, s36_1_1, s36_2_2, c36_2_2);
	full_adder ad36_2_3(s36_1_2, s36_1_3, s36_1_4, s36_2_3, c36_2_3);
	full_adder ad37_2_0(c36_1_0, c36_1_1, c36_1_2, s37_2_0, c37_2_0);
	full_adder ad37_2_1(c36_1_3, c36_1_4, c36_1_5, s37_2_1, c37_2_1);
	full_adder ad37_2_2(s37_1_0, s37_1_1, s37_1_2, s37_2_2, c37_2_2);
	full_adder ad37_2_3(s37_1_3, s37_1_4, s37_1_5, s37_2_3, c37_2_3);
	full_adder ad38_2_0(c37_1_0, c37_1_1, c37_1_2, s38_2_0, c38_2_0);
	full_adder ad38_2_1(c37_1_3, c37_1_4, c37_1_5, s38_2_1, c38_2_1);
	full_adder ad38_2_2(s38_1_0, s38_1_1, s38_1_2, s38_2_2, c38_2_2);
	full_adder ad38_2_3(s38_1_3, s38_1_4, s38_1_5, s38_2_3, c38_2_3);
	full_adder ad39_2_0(c38_1_0, c38_1_1, c38_1_2, s39_2_0, c39_2_0);
	full_adder ad39_2_1(c38_1_3, c38_1_4, c38_1_5, s39_2_1, c39_2_1);
	full_adder ad39_2_2(s39_1_0, s39_1_1, s39_1_2, s39_2_2, c39_2_2);
	full_adder ad39_2_3(s39_1_3, s39_1_4, s39_0_7, s39_2_3, c39_2_3);
	full_adder ad40_2_0(c39_1_0, c39_1_1, c39_1_2, s40_2_0, c40_2_0);
	full_adder ad40_2_1(c39_1_3, c39_1_4, s40_1_0, s40_2_1, c40_2_1);
	full_adder ad40_2_2(s40_1_1, s40_1_2, s40_1_3, s40_2_2, c40_2_2);
	half_adder ha40_2_3(s40_1_4, s40_0_7, s40_2_3, c40_2_3);
	full_adder ad41_2_0(c40_1_0, c40_1_1, c40_1_2, s41_2_0, c41_2_0);
	full_adder ad41_2_1(c40_1_3, c40_1_4, s41_1_0, s41_2_1, c41_2_1);
	full_adder ad41_2_2(s41_1_1, s41_1_2, s41_1_3, s41_2_2, c41_2_2);
	half_adder ha41_2_3(s41_1_4, a31_41, s41_2_3, c41_2_3);
	full_adder ad42_2_0(c41_1_0, c41_1_1, c41_1_2, s42_2_0, c42_2_0);
	full_adder ad42_2_1(c41_1_3, c41_1_4, s42_1_0, s42_2_1, c42_2_1);
	full_adder ad42_2_2(s42_1_1, s42_1_2, s42_1_3, s42_2_2, c42_2_2);
	full_adder ad43_2_0(c42_1_0, c42_1_1, c42_1_2, s43_2_0, c43_2_0);
	full_adder ad43_2_1(c42_1_3, c42_1_4, s43_1_0, s43_2_1, c43_2_1);
	full_adder ad43_2_2(s43_1_1, s43_1_2, s43_1_3, s43_2_2, c43_2_2);
	full_adder ad44_2_0(c43_1_0, c43_1_1, c43_1_2, s44_2_0, c44_2_0);
	full_adder ad44_2_1(c43_1_3, c43_1_4, s44_1_0, s44_2_1, c44_2_1);
	full_adder ad44_2_2(s44_1_1, s44_1_2, s44_1_3, s44_2_2, c44_2_2);
	full_adder ad45_2_0(c44_1_0, c44_1_1, c44_1_2, s45_2_0, c45_2_0);
	full_adder ad45_2_1(c44_1_3, c44_1_4, s45_1_0, s45_2_1, c45_2_1);
	full_adder ad45_2_2(s45_1_1, s45_1_2, s45_1_3, s45_2_2, c45_2_2);
	full_adder ad46_2_0(c45_1_0, c45_1_1, c45_1_2, s46_2_0, c46_2_0);
	full_adder ad46_2_1(c45_1_3, s46_1_0, s46_1_1, s46_2_1, c46_2_1);
	half_adder ha46_2_2(s46_1_2, s46_1_3, s46_2_2, c46_2_2);
	full_adder ad47_2_0(c46_1_0, c46_1_1, c46_1_2, s47_2_0, c47_2_0);
	full_adder ad47_2_1(c46_1_3, s47_1_0, s47_1_1, s47_2_1, c47_2_1);
	half_adder ha47_2_2(s47_1_2, s47_1_3, s47_2_2, c47_2_2);
	full_adder ad48_2_0(c47_1_0, c47_1_1, c47_1_2, s48_2_0, c48_2_0);
	full_adder ad48_2_1(c47_1_3, s48_1_0, s48_1_1, s48_2_1, c48_2_1);
	half_adder ha48_2_2(s48_1_2, s48_0_4, s48_2_2, c48_2_2);
	full_adder ad49_2_0(c48_1_0, c48_1_1, c48_1_2, s49_2_0, c49_2_0);
	full_adder ad49_2_1(s49_1_0, s49_1_1, s49_1_2, s49_2_1, c49_2_1);
	full_adder ad50_2_0(c49_1_0, c49_1_1, c49_1_2, s50_2_0, c50_2_0);
	full_adder ad50_2_1(s50_1_0, s50_1_1, s50_1_2, s50_2_1, c50_2_1);
	full_adder ad51_2_0(c50_1_0, c50_1_1, c50_1_2, s51_2_0, c51_2_0);
	full_adder ad51_2_1(s51_1_0, s51_1_1, s51_1_2, s51_2_1, c51_2_1);
	full_adder ad52_2_0(c51_1_0, c51_1_1, c51_1_2, s52_2_0, c52_2_0);
	full_adder ad52_2_1(s52_1_0, s52_1_1, s52_1_2, s52_2_1, c52_2_1);
	full_adder ad53_2_0(c52_1_0, c52_1_1, c52_1_2, s53_2_0, c53_2_0);
	full_adder ad53_2_1(s53_1_0, s53_1_1, s53_1_2, s53_2_1, c53_2_1);
	full_adder ad54_2_0(c53_1_0, c53_1_1, c53_1_2, s54_2_0, c54_2_0);
	half_adder ha54_2_1(s54_1_0, s54_1_1, s54_2_1, c54_2_1);
	full_adder ad55_2_0(c54_1_0, c54_1_1, s55_1_0, s55_2_0, c55_2_0);
	full_adder ad56_2_0(c55_1_0, c55_1_1, s56_1_0, s56_2_0, c56_2_0);
	full_adder ad57_2_0(c56_1_0, c56_1_1, s57_1_0, s57_2_0, c57_2_0);
	full_adder ad58_2_0(c57_1_0, s58_1_0, s58_0_1, s58_2_0, c58_2_0);
	full_adder ad59_2_0(c58_1_0, s59_1_0, a31_59, s59_2_0, c59_2_0);
	half_adder ha60_2_0(c59_1_0, s60_1_0, s60_2_0, c60_2_0);
	half_adder ha61_2_0(c60_1_0, s61_1_0, s61_2_0, c61_2_0);
	half_adder ha62_2_0(c61_1_0, s62_1_0, s62_2_0, c62_2_0);
	half_adder ha63_2_0(c62_1_0, 1'b1, s63_2_0, c63_2_0);

	half_adder ha4_3_0(c3_2_0, s4_2_0, s4_3_0, c4_3_0);
	half_adder ha5_3_0(c4_2_0, s5_2_0, s5_3_0, c5_3_0);
	half_adder ha6_3_0(c5_2_0, s6_2_0, s6_3_0, c6_3_0);
	full_adder ad7_3_0(c6_2_0, s7_2_0, s7_1_1, s7_3_0, c7_3_0);
	full_adder ad8_3_0(c7_2_0, s8_2_0, s8_1_1, s8_3_0, c8_3_0);
	full_adder ad9_3_0(c8_2_0, s9_2_0, s9_2_1, s9_3_0, c9_3_0);
	full_adder ad10_3_0(c9_2_0, c9_2_1, s10_2_0, s10_3_0, c10_3_0);
	full_adder ad11_3_0(c10_2_0, c10_2_1, s11_2_0, s11_3_0, c11_3_0);
	full_adder ad12_3_0(c11_2_0, c11_2_1, s12_2_0, s12_3_0, c12_3_0);
	full_adder ad13_3_0(c12_2_0, c12_2_1, s13_2_0, s13_3_0, c13_3_0);
	full_adder ad14_3_0(c13_2_0, c13_2_1, s14_2_0, s14_3_0, c14_3_0);
	half_adder ha14_3_1(s14_2_1, s14_0_4, s14_3_1, c14_3_1);
	full_adder ad15_3_0(c14_2_0, c14_2_1, s15_2_0, s15_3_0, c15_3_0);
	half_adder ha15_3_1(s15_2_1, s15_1_3, s15_3_1, c15_3_1);
	full_adder ad16_3_0(c15_2_0, c15_2_1, s16_2_0, s16_3_0, c16_3_0);
	half_adder ha16_3_1(s16_2_1, s16_2_2, s16_3_1, c16_3_1);
	full_adder ad17_3_0(c16_2_0, c16_2_1, c16_2_2, s17_3_0, c17_3_0);
	full_adder ad17_3_1(s17_2_0, s17_2_1, s17_2_2, s17_3_1, c17_3_1);
	full_adder ad18_3_0(c17_2_0, c17_2_1, c17_2_2, s18_3_0, c18_3_0);
	full_adder ad18_3_1(s18_2_0, s18_2_1, s18_2_2, s18_3_1, c18_3_1);
	full_adder ad19_3_0(c18_2_0, c18_2_1, c18_2_2, s19_3_0, c19_3_0);
	full_adder ad19_3_1(s19_2_0, s19_2_1, s19_2_2, s19_3_1, c19_3_1);
	full_adder ad20_3_0(c19_2_0, c19_2_1, c19_2_2, s20_3_0, c20_3_0);
	full_adder ad20_3_1(s20_2_0, s20_2_1, s20_2_2, s20_3_1, c20_3_1);
	full_adder ad21_3_0(c20_2_0, c20_2_1, c20_2_2, s21_3_0, c21_3_0);
	full_adder ad21_3_1(s21_2_0, s21_2_1, s21_2_2, s21_3_1, c21_3_1);
	full_adder ad22_3_0(c21_2_0, c21_2_1, c21_2_2, s22_3_0, c22_3_0);
	full_adder ad22_3_1(s22_2_0, s22_2_1, s22_2_2, s22_3_1, c22_3_1);
	full_adder ad23_3_0(c22_2_0, c22_2_1, c22_2_2, s23_3_0, c23_3_0);
	full_adder ad23_3_1(s23_2_0, s23_2_1, s23_2_2, s23_3_1, c23_3_1);
	full_adder ad24_3_0(c23_2_0, c23_2_1, c23_2_2, s24_3_0, c24_3_0);
	full_adder ad24_3_1(c23_2_3, s24_2_0, s24_2_1, s24_3_1, c24_3_1);
	half_adder ha24_3_2(s24_2_2, s24_2_3, s24_3_2, c24_3_2);
	full_adder ad25_3_0(c24_2_0, c24_2_1, c24_2_2, s25_3_0, c25_3_0);
	full_adder ad25_3_1(c24_2_3, s25_2_0, s25_2_1, s25_3_1, c25_3_1);
	half_adder ha25_3_2(s25_2_2, s25_2_3, s25_3_2, c25_3_2);
	full_adder ad26_3_0(c25_2_0, c25_2_1, c25_2_2, s26_3_0, c26_3_0);
	full_adder ad26_3_1(c25_2_3, s26_2_0, s26_2_1, s26_3_1, c26_3_1);
	half_adder ha26_3_2(s26_2_2, s26_2_3, s26_3_2, c26_3_2);
	full_adder ad27_3_0(c26_2_0, c26_2_1, c26_2_2, s27_3_0, c27_3_0);
	full_adder ad27_3_1(c26_2_3, s27_2_0, s27_2_1, s27_3_1, c27_3_1);
	full_adder ad27_3_2(s27_2_2, s27_2_3, a27_27, s27_3_2, c27_3_2);
	full_adder ad28_3_0(c27_2_0, c27_2_1, c27_2_2, s28_3_0, c28_3_0);
	full_adder ad28_3_1(c27_2_3, s28_2_0, s28_2_1, s28_3_1, c28_3_1);
	full_adder ad28_3_2(s28_2_2, s28_2_3, s28_0_9, s28_3_2, c28_3_2);
	full_adder ad29_3_0(c28_2_0, c28_2_1, c28_2_2, s29_3_0, c29_3_0);
	full_adder ad29_3_1(c28_2_3, s29_2_0, s29_2_1, s29_3_1, c29_3_1);
	full_adder ad29_3_2(s29_2_2, s29_2_3, s29_1_6, s29_3_2, c29_3_2);
	full_adder ad30_3_0(c29_2_0, c29_2_1, c29_2_2, s30_3_0, c30_3_0);
	full_adder ad30_3_1(c29_2_3, s30_2_0, s30_2_1, s30_3_1, c30_3_1);
	full_adder ad30_3_2(s30_2_2, s30_2_3, s30_2_4, s30_3_2, c30_3_2);
	full_adder ad31_3_0(c30_2_0, c30_2_1, c30_2_2, s31_3_0, c31_3_0);
	full_adder ad31_3_1(c30_2_3, c30_2_4, s31_2_0, s31_3_1, c31_3_1);
	full_adder ad31_3_2(s31_2_1, s31_2_2, s31_2_3, s31_3_2, c31_3_2);
	full_adder ad32_3_0(c31_2_0, c31_2_1, c31_2_2, s32_3_0, c32_3_0);
	full_adder ad32_3_1(c31_2_3, c31_2_4, s32_2_0, s32_3_1, c32_3_1);
	full_adder ad32_3_2(s32_2_1, s32_2_2, s32_2_3, s32_3_2, c32_3_2);
	full_adder ad33_3_0(c32_2_0, c32_2_1, c32_2_2, s33_3_0, c33_3_0);
	full_adder ad33_3_1(c32_2_3, c32_2_4, s33_2_0, s33_3_1, c33_3_1);
	full_adder ad33_3_2(s33_2_1, s33_2_2, s33_2_3, s33_3_2, c33_3_2);
	full_adder ad34_3_0(c33_2_0, c33_2_1, c33_2_2, s34_3_0, c34_3_0);
	full_adder ad34_3_1(c33_2_3, c33_2_4, s34_2_0, s34_3_1, c34_3_1);
	full_adder ad34_3_2(s34_2_1, s34_2_2, s34_2_3, s34_3_2, c34_3_2);
	full_adder ad35_3_0(c34_2_0, c34_2_1, c34_2_2, s35_3_0, c35_3_0);
	full_adder ad35_3_1(c34_2_3, c34_2_4, s35_2_0, s35_3_1, c35_3_1);
	full_adder ad35_3_2(s35_2_1, s35_2_2, s35_2_3, s35_3_2, c35_3_2);
	full_adder ad36_3_0(c35_2_0, c35_2_1, c35_2_2, s36_3_0, c36_3_0);
	full_adder ad36_3_1(c35_2_3, c35_2_4, s36_2_0, s36_3_1, c36_3_1);
	full_adder ad36_3_2(s36_2_1, s36_2_2, s36_2_3, s36_3_2, c36_3_2);
	full_adder ad37_3_0(c36_2_0, c36_2_1, c36_2_2, s37_3_0, c37_3_0);
	full_adder ad37_3_1(c36_2_3, s37_2_0, s37_2_1, s37_3_1, c37_3_1);
	half_adder ha37_3_2(s37_2_2, s37_2_3, s37_3_2, c37_3_2);
	full_adder ad38_3_0(c37_2_0, c37_2_1, c37_2_2, s38_3_0, c38_3_0);
	full_adder ad38_3_1(c37_2_3, s38_2_0, s38_2_1, s38_3_1, c38_3_1);
	half_adder ha38_3_2(s38_2_2, s38_2_3, s38_3_2, c38_3_2);
	full_adder ad39_3_0(c38_2_0, c38_2_1, c38_2_2, s39_3_0, c39_3_0);
	full_adder ad39_3_1(c38_2_3, s39_2_0, s39_2_1, s39_3_1, c39_3_1);
	half_adder ha39_3_2(s39_2_2, s39_2_3, s39_3_2, c39_3_2);
	full_adder ad40_3_0(c39_2_0, c39_2_1, c39_2_2, s40_3_0, c40_3_0);
	full_adder ad40_3_1(c39_2_3, s40_2_0, s40_2_1, s40_3_1, c40_3_1);
	half_adder ha40_3_2(s40_2_2, s40_2_3, s40_3_2, c40_3_2);
	full_adder ad41_3_0(c40_2_0, c40_2_1, c40_2_2, s41_3_0, c41_3_0);
	full_adder ad41_3_1(c40_2_3, s41_2_0, s41_2_1, s41_3_1, c41_3_1);
	half_adder ha41_3_2(s41_2_2, s41_2_3, s41_3_2, c41_3_2);
	full_adder ad42_3_0(c41_2_0, c41_2_1, c41_2_2, s42_3_0, c42_3_0);
	full_adder ad42_3_1(c41_2_3, s42_2_0, s42_2_1, s42_3_1, c42_3_1);
	half_adder ha42_3_2(s42_2_2, s42_1_4, s42_3_2, c42_3_2);
	full_adder ad43_3_0(c42_2_0, c42_2_1, c42_2_2, s43_3_0, c43_3_0);
	full_adder ad43_3_1(s43_2_0, s43_2_1, s43_2_2, s43_3_1, c43_3_1);
	full_adder ad44_3_0(c43_2_0, c43_2_1, c43_2_2, s44_3_0, c44_3_0);
	full_adder ad44_3_1(s44_2_0, s44_2_1, s44_2_2, s44_3_1, c44_3_1);
	full_adder ad45_3_0(c44_2_0, c44_2_1, c44_2_2, s45_3_0, c45_3_0);
	full_adder ad45_3_1(s45_2_0, s45_2_1, s45_2_2, s45_3_1, c45_3_1);
	full_adder ad46_3_0(c45_2_0, c45_2_1, c45_2_2, s46_3_0, c46_3_0);
	full_adder ad46_3_1(s46_2_0, s46_2_1, s46_2_2, s46_3_1, c46_3_1);
	full_adder ad47_3_0(c46_2_0, c46_2_1, c46_2_2, s47_3_0, c47_3_0);
	full_adder ad47_3_1(s47_2_0, s47_2_1, s47_2_2, s47_3_1, c47_3_1);
	full_adder ad48_3_0(c47_2_0, c47_2_1, c47_2_2, s48_3_0, c48_3_0);
	full_adder ad48_3_1(s48_2_0, s48_2_1, s48_2_2, s48_3_1, c48_3_1);
	full_adder ad49_3_0(c48_2_0, c48_2_1, c48_2_2, s49_3_0, c49_3_0);
	full_adder ad49_3_1(s49_2_0, s49_2_1, s49_0_4, s49_3_1, c49_3_1);
	full_adder ad50_3_0(c49_2_0, c49_2_1, s50_2_0, s50_3_0, c50_3_0);
	half_adder ha50_3_1(s50_2_1, a31_50, s50_3_1, c50_3_1);
	full_adder ad51_3_0(c50_2_0, c50_2_1, s51_2_0, s51_3_0, c51_3_0);
	full_adder ad52_3_0(c51_2_0, c51_2_1, s52_2_0, s52_3_0, c52_3_0);
	full_adder ad53_3_0(c52_2_0, c52_2_1, s53_2_0, s53_3_0, c53_3_0);
	full_adder ad54_3_0(c53_2_0, c53_2_1, s54_2_0, s54_3_0, c54_3_0);
	full_adder ad55_3_0(c54_2_0, c54_2_1, s55_2_0, s55_3_0, c55_3_0);
	full_adder ad56_3_0(c55_2_0, s56_2_0, s56_1_1, s56_3_0, c56_3_0);
	full_adder ad57_3_0(c56_2_0, s57_2_0, s57_0_1, s57_3_0, c57_3_0);
	half_adder ha58_3_0(c57_2_0, s58_2_0, s58_3_0, c58_3_0);
	half_adder ha59_3_0(c58_2_0, s59_2_0, s59_3_0, c59_3_0);
	half_adder ha60_3_0(c59_2_0, s60_2_0, s60_3_0, c60_3_0);
	half_adder ha61_3_0(c60_2_0, s61_2_0, s61_3_0, c61_3_0);
	half_adder ha62_3_0(c61_2_0, s62_2_0, s62_3_0, c62_3_0);
	half_adder ha63_3_0(c62_2_0, s63_2_0, s63_3_0, c63_3_0);

	half_adder ha5_4_0(c4_3_0, s5_3_0, s5_4_0, c5_4_0);
	half_adder ha6_4_0(c5_3_0, s6_3_0, s6_4_0, c6_4_0);
	half_adder ha7_4_0(c6_3_0, s7_3_0, s7_4_0, c7_4_0);
	half_adder ha8_4_0(c7_3_0, s8_3_0, s8_4_0, c8_4_0);
	half_adder ha9_4_0(c8_3_0, s9_3_0, s9_4_0, c9_4_0);
	full_adder ad10_4_0(c9_3_0, s10_3_0, s10_2_1, s10_4_0, c10_4_0);
	full_adder ad11_4_0(c10_3_0, s11_3_0, s11_2_1, s11_4_0, c11_4_0);
	full_adder ad12_4_0(c11_3_0, s12_3_0, s12_2_1, s12_4_0, c12_4_0);
	full_adder ad13_4_0(c12_3_0, s13_3_0, s13_2_1, s13_4_0, c13_4_0);
	full_adder ad14_4_0(c13_3_0, s14_3_0, s14_3_1, s14_4_0, c14_4_0);
	full_adder ad15_4_0(c14_3_0, c14_3_1, s15_3_0, s15_4_0, c15_4_0);
	full_adder ad16_4_0(c15_3_0, c15_3_1, s16_3_0, s16_4_0, c16_4_0);
	full_adder ad17_4_0(c16_3_0, c16_3_1, s17_3_0, s17_4_0, c17_4_0);
	full_adder ad18_4_0(c17_3_0, c17_3_1, s18_3_0, s18_4_0, c18_4_0);
	full_adder ad19_4_0(c18_3_0, c18_3_1, s19_3_0, s19_4_0, c19_4_0);
	full_adder ad20_4_0(c19_3_0, c19_3_1, s20_3_0, s20_4_0, c20_4_0);
	full_adder ad21_4_0(c20_3_0, c20_3_1, s21_3_0, s21_4_0, c21_4_0);
	half_adder ha21_4_1(s21_3_1, s21_1_4, s21_4_1, c21_4_1);
	full_adder ad22_4_0(c21_3_0, c21_3_1, s22_3_0, s22_4_0, c22_4_0);
	half_adder ha22_4_1(s22_3_1, s22_1_4, s22_4_1, c22_4_1);
	full_adder ad23_4_0(c22_3_0, c22_3_1, s23_3_0, s23_4_0, c23_4_0);
	half_adder ha23_4_1(s23_3_1, s23_2_3, s23_4_1, c23_4_1);
	full_adder ad24_4_0(c23_3_0, c23_3_1, s24_3_0, s24_4_0, c24_4_0);
	half_adder ha24_4_1(s24_3_1, s24_3_2, s24_4_1, c24_4_1);
	full_adder ad25_4_0(c24_3_0, c24_3_1, c24_3_2, s25_4_0, c25_4_0);
	full_adder ad25_4_1(s25_3_0, s25_3_1, s25_3_2, s25_4_1, c25_4_1);
	full_adder ad26_4_0(c25_3_0, c25_3_1, c25_3_2, s26_4_0, c26_4_0);
	full_adder ad26_4_1(s26_3_0, s26_3_1, s26_3_2, s26_4_1, c26_4_1);
	full_adder ad27_4_0(c26_3_0, c26_3_1, c26_3_2, s27_4_0, c27_4_0);
	full_adder ad27_4_1(s27_3_0, s27_3_1, s27_3_2, s27_4_1, c27_4_1);
	full_adder ad28_4_0(c27_3_0, c27_3_1, c27_3_2, s28_4_0, c28_4_0);
	full_adder ad28_4_1(s28_3_0, s28_3_1, s28_3_2, s28_4_1, c28_4_1);
	full_adder ad29_4_0(c28_3_0, c28_3_1, c28_3_2, s29_4_0, c29_4_0);
	full_adder ad29_4_1(s29_3_0, s29_3_1, s29_3_2, s29_4_1, c29_4_1);
	full_adder ad30_4_0(c29_3_0, c29_3_1, c29_3_2, s30_4_0, c30_4_0);
	full_adder ad30_4_1(s30_3_0, s30_3_1, s30_3_2, s30_4_1, c30_4_1);
	full_adder ad31_4_0(c30_3_0, c30_3_1, c30_3_2, s31_4_0, c31_4_0);
	full_adder ad31_4_1(s31_3_0, s31_3_1, s31_3_2, s31_4_1, c31_4_1);
	full_adder ad32_4_0(c31_3_0, c31_3_1, c31_3_2, s32_4_0, c32_4_0);
	full_adder ad32_4_1(s32_3_0, s32_3_1, s32_3_2, s32_4_1, c32_4_1);
	full_adder ad33_4_0(c32_3_0, c32_3_1, c32_3_2, s33_4_0, c33_4_0);
	full_adder ad33_4_1(s33_3_0, s33_3_1, s33_3_2, s33_4_1, c33_4_1);
	full_adder ad34_4_0(c33_3_0, c33_3_1, c33_3_2, s34_4_0, c34_4_0);
	full_adder ad34_4_1(s34_3_0, s34_3_1, s34_3_2, s34_4_1, c34_4_1);
	full_adder ad35_4_0(c34_3_0, c34_3_1, c34_3_2, s35_4_0, c35_4_0);
	full_adder ad35_4_1(s35_3_0, s35_3_1, s35_3_2, s35_4_1, c35_4_1);
	full_adder ad36_4_0(c35_3_0, c35_3_1, c35_3_2, s36_4_0, c36_4_0);
	full_adder ad36_4_1(s36_3_0, s36_3_1, s36_3_2, s36_4_1, c36_4_1);
	full_adder ad37_4_0(c36_3_0, c36_3_1, c36_3_2, s37_4_0, c37_4_0);
	full_adder ad37_4_1(s37_3_0, s37_3_1, s37_3_2, s37_4_1, c37_4_1);
	full_adder ad38_4_0(c37_3_0, c37_3_1, c37_3_2, s38_4_0, c38_4_0);
	full_adder ad38_4_1(s38_3_0, s38_3_1, s38_3_2, s38_4_1, c38_4_1);
	full_adder ad39_4_0(c38_3_0, c38_3_1, c38_3_2, s39_4_0, c39_4_0);
	full_adder ad39_4_1(s39_3_0, s39_3_1, s39_3_2, s39_4_1, c39_4_1);
	full_adder ad40_4_0(c39_3_0, c39_3_1, c39_3_2, s40_4_0, c40_4_0);
	full_adder ad40_4_1(s40_3_0, s40_3_1, s40_3_2, s40_4_1, c40_4_1);
	full_adder ad41_4_0(c40_3_0, c40_3_1, c40_3_2, s41_4_0, c41_4_0);
	full_adder ad41_4_1(s41_3_0, s41_3_1, s41_3_2, s41_4_1, c41_4_1);
	full_adder ad42_4_0(c41_3_0, c41_3_1, c41_3_2, s42_4_0, c42_4_0);
	full_adder ad42_4_1(s42_3_0, s42_3_1, s42_3_2, s42_4_1, c42_4_1);
	full_adder ad43_4_0(c42_3_0, c42_3_1, c42_3_2, s43_4_0, c43_4_0);
	full_adder ad43_4_1(s43_3_0, s43_3_1, s43_1_4, s43_4_1, c43_4_1);
	full_adder ad44_4_0(c43_3_0, c43_3_1, s44_3_0, s44_4_0, c44_4_0);
	half_adder ha44_4_1(s44_3_1, s44_1_4, s44_4_1, c44_4_1);
	full_adder ad45_4_0(c44_3_0, c44_3_1, s45_3_0, s45_4_0, c45_4_0);
	full_adder ad46_4_0(c45_3_0, c45_3_1, s46_3_0, s46_4_0, c46_4_0);
	full_adder ad47_4_0(c46_3_0, c46_3_1, s47_3_0, s47_4_0, c47_4_0);
	full_adder ad48_4_0(c47_3_0, c47_3_1, s48_3_0, s48_4_0, c48_4_0);
	full_adder ad49_4_0(c48_3_0, c48_3_1, s49_3_0, s49_4_0, c49_4_0);
	full_adder ad50_4_0(c49_3_0, c49_3_1, s50_3_0, s50_4_0, c50_4_0);
	full_adder ad51_4_0(c50_3_0, c50_3_1, s51_3_0, s51_4_0, c51_4_0);
	full_adder ad52_4_0(c51_3_0, s52_3_0, s52_2_1, s52_4_0, c52_4_0);
	full_adder ad53_4_0(c52_3_0, s53_3_0, s53_2_1, s53_4_0, c53_4_0);
	full_adder ad54_4_0(c53_3_0, s54_3_0, s54_2_1, s54_4_0, c54_4_0);
	full_adder ad55_4_0(c54_3_0, s55_3_0, s55_1_1, s55_4_0, c55_4_0);
	half_adder ha56_4_0(c55_3_0, s56_3_0, s56_4_0, c56_4_0);
	half_adder ha57_4_0(c56_3_0, s57_3_0, s57_4_0, c57_4_0);
	half_adder ha58_4_0(c57_3_0, s58_3_0, s58_4_0, c58_4_0);
	half_adder ha59_4_0(c58_3_0, s59_3_0, s59_4_0, c59_4_0);
	half_adder ha60_4_0(c59_3_0, s60_3_0, s60_4_0, c60_4_0);
	half_adder ha61_4_0(c60_3_0, s61_3_0, s61_4_0, c61_4_0);
	half_adder ha62_4_0(c61_3_0, s62_3_0, s62_4_0, c62_4_0);
	half_adder ha63_4_0(c62_3_0, s63_3_0, s63_4_0, c63_4_0);

	half_adder ha6_5_0(c5_4_0, s6_4_0, s6_5_0, c6_5_0);
	half_adder ha7_5_0(c6_4_0, s7_4_0, s7_5_0, c7_5_0);
	half_adder ha8_5_0(c7_4_0, s8_4_0, s8_5_0, c8_5_0);
	half_adder ha9_5_0(c8_4_0, s9_4_0, s9_5_0, c9_5_0);
	half_adder ha10_5_0(c9_4_0, s10_4_0, s10_5_0, c10_5_0);
	half_adder ha11_5_0(c10_4_0, s11_4_0, s11_5_0, c11_5_0);
	half_adder ha12_5_0(c11_4_0, s12_4_0, s12_5_0, c12_5_0);
	half_adder ha13_5_0(c12_4_0, s13_4_0, s13_5_0, c13_5_0);
	half_adder ha14_5_0(c13_4_0, s14_4_0, s14_5_0, c14_5_0);
	full_adder ad15_5_0(c14_4_0, s15_4_0, s15_3_1, s15_5_0, c15_5_0);
	full_adder ad16_5_0(c15_4_0, s16_4_0, s16_3_1, s16_5_0, c16_5_0);
	full_adder ad17_5_0(c16_4_0, s17_4_0, s17_3_1, s17_5_0, c17_5_0);
	full_adder ad18_5_0(c17_4_0, s18_4_0, s18_3_1, s18_5_0, c18_5_0);
	full_adder ad19_5_0(c18_4_0, s19_4_0, s19_3_1, s19_5_0, c19_5_0);
	full_adder ad20_5_0(c19_4_0, s20_4_0, s20_3_1, s20_5_0, c20_5_0);
	full_adder ad21_5_0(c20_4_0, s21_4_0, s21_4_1, s21_5_0, c21_5_0);
	full_adder ad22_5_0(c21_4_0, c21_4_1, s22_4_0, s22_5_0, c22_5_0);
	full_adder ad23_5_0(c22_4_0, c22_4_1, s23_4_0, s23_5_0, c23_5_0);
	full_adder ad24_5_0(c23_4_0, c23_4_1, s24_4_0, s24_5_0, c24_5_0);
	full_adder ad25_5_0(c24_4_0, c24_4_1, s25_4_0, s25_5_0, c25_5_0);
	full_adder ad26_5_0(c25_4_0, c25_4_1, s26_4_0, s26_5_0, c26_5_0);
	full_adder ad27_5_0(c26_4_0, c26_4_1, s27_4_0, s27_5_0, c27_5_0);
	full_adder ad28_5_0(c27_4_0, c27_4_1, s28_4_0, s28_5_0, c28_5_0);
	full_adder ad29_5_0(c28_4_0, c28_4_1, s29_4_0, s29_5_0, c29_5_0);
	full_adder ad30_5_0(c29_4_0, c29_4_1, s30_4_0, s30_5_0, c30_5_0);
	full_adder ad31_5_0(c30_4_0, c30_4_1, s31_4_0, s31_5_0, c31_5_0);
	half_adder ha31_5_1(s31_4_1, s31_2_4, s31_5_1, c31_5_1);
	full_adder ad32_5_0(c31_4_0, c31_4_1, s32_4_0, s32_5_0, c32_5_0);
	half_adder ha32_5_1(s32_4_1, s32_2_4, s32_5_1, c32_5_1);
	full_adder ad33_5_0(c32_4_0, c32_4_1, s33_4_0, s33_5_0, c33_5_0);
	half_adder ha33_5_1(s33_4_1, s33_2_4, s33_5_1, c33_5_1);
	full_adder ad34_5_0(c33_4_0, c33_4_1, s34_4_0, s34_5_0, c34_5_0);
	half_adder ha34_5_1(s34_4_1, s34_2_4, s34_5_1, c34_5_1);
	full_adder ad35_5_0(c34_4_0, c34_4_1, s35_4_0, s35_5_0, c35_5_0);
	half_adder ha35_5_1(s35_4_1, s35_2_4, s35_5_1, c35_5_1);
	full_adder ad36_5_0(c35_4_0, c35_4_1, s36_4_0, s36_5_0, c36_5_0);
	half_adder ha36_5_1(s36_4_1, s36_1_5, s36_5_1, c36_5_1);
	full_adder ad37_5_0(c36_4_0, c36_4_1, s37_4_0, s37_5_0, c37_5_0);
	full_adder ad38_5_0(c37_4_0, c37_4_1, s38_4_0, s38_5_0, c38_5_0);
	full_adder ad39_5_0(c38_4_0, c38_4_1, s39_4_0, s39_5_0, c39_5_0);
	full_adder ad40_5_0(c39_4_0, c39_4_1, s40_4_0, s40_5_0, c40_5_0);
	full_adder ad41_5_0(c40_4_0, c40_4_1, s41_4_0, s41_5_0, c41_5_0);
	full_adder ad42_5_0(c41_4_0, c41_4_1, s42_4_0, s42_5_0, c42_5_0);
	full_adder ad43_5_0(c42_4_0, c42_4_1, s43_4_0, s43_5_0, c43_5_0);
	full_adder ad44_5_0(c43_4_0, c43_4_1, s44_4_0, s44_5_0, c44_5_0);
	full_adder ad45_5_0(c44_4_0, c44_4_1, s45_4_0, s45_5_0, c45_5_0);
	full_adder ad46_5_0(c45_4_0, s46_4_0, s46_3_1, s46_5_0, c46_5_0);
	full_adder ad47_5_0(c46_4_0, s47_4_0, s47_3_1, s47_5_0, c47_5_0);
	full_adder ad48_5_0(c47_4_0, s48_4_0, s48_3_1, s48_5_0, c48_5_0);
	full_adder ad49_5_0(c48_4_0, s49_4_0, s49_3_1, s49_5_0, c49_5_0);
	full_adder ad50_5_0(c49_4_0, s50_4_0, s50_3_1, s50_5_0, c50_5_0);
	full_adder ad51_5_0(c50_4_0, s51_4_0, s51_2_1, s51_5_0, c51_5_0);
	half_adder ha52_5_0(c51_4_0, s52_4_0, s52_5_0, c52_5_0);
	half_adder ha53_5_0(c52_4_0, s53_4_0, s53_5_0, c53_5_0);
	half_adder ha54_5_0(c53_4_0, s54_4_0, s54_5_0, c54_5_0);
	half_adder ha55_5_0(c54_4_0, s55_4_0, s55_5_0, c55_5_0);
	half_adder ha56_5_0(c55_4_0, s56_4_0, s56_5_0, c56_5_0);
	half_adder ha57_5_0(c56_4_0, s57_4_0, s57_5_0, c57_5_0);
	half_adder ha58_5_0(c57_4_0, s58_4_0, s58_5_0, c58_5_0);
	half_adder ha59_5_0(c58_4_0, s59_4_0, s59_5_0, c59_5_0);
	half_adder ha60_5_0(c59_4_0, s60_4_0, s60_5_0, c60_5_0);
	half_adder ha61_5_0(c60_4_0, s61_4_0, s61_5_0, c61_5_0);
	half_adder ha62_5_0(c61_4_0, s62_4_0, s62_5_0, c62_5_0);
	half_adder ha63_5_0(c62_4_0, s63_4_0, s63_5_0, c63_5_0);

	half_adder ha7_6_0(c6_5_0, s7_5_0, s7_6_0, c7_6_0);
	half_adder ha8_6_0(c7_5_0, s8_5_0, s8_6_0, c8_6_0);
	half_adder ha9_6_0(c8_5_0, s9_5_0, s9_6_0, c9_6_0);
	half_adder ha10_6_0(c9_5_0, s10_5_0, s10_6_0, c10_6_0);
	half_adder ha11_6_0(c10_5_0, s11_5_0, s11_6_0, c11_6_0);
	half_adder ha12_6_0(c11_5_0, s12_5_0, s12_6_0, c12_6_0);
	half_adder ha13_6_0(c12_5_0, s13_5_0, s13_6_0, c13_6_0);
	half_adder ha14_6_0(c13_5_0, s14_5_0, s14_6_0, c14_6_0);
	half_adder ha15_6_0(c14_5_0, s15_5_0, s15_6_0, c15_6_0);
	half_adder ha16_6_0(c15_5_0, s16_5_0, s16_6_0, c16_6_0);
	half_adder ha17_6_0(c16_5_0, s17_5_0, s17_6_0, c17_6_0);
	half_adder ha18_6_0(c17_5_0, s18_5_0, s18_6_0, c18_6_0);
	half_adder ha19_6_0(c18_5_0, s19_5_0, s19_6_0, c19_6_0);
	half_adder ha20_6_0(c19_5_0, s20_5_0, s20_6_0, c20_6_0);
	half_adder ha21_6_0(c20_5_0, s21_5_0, s21_6_0, c21_6_0);
	full_adder ad22_6_0(c21_5_0, s22_5_0, s22_4_1, s22_6_0, c22_6_0);
	full_adder ad23_6_0(c22_5_0, s23_5_0, s23_4_1, s23_6_0, c23_6_0);
	full_adder ad24_6_0(c23_5_0, s24_5_0, s24_4_1, s24_6_0, c24_6_0);
	full_adder ad25_6_0(c24_5_0, s25_5_0, s25_4_1, s25_6_0, c25_6_0);
	full_adder ad26_6_0(c25_5_0, s26_5_0, s26_4_1, s26_6_0, c26_6_0);
	full_adder ad27_6_0(c26_5_0, s27_5_0, s27_4_1, s27_6_0, c27_6_0);
	full_adder ad28_6_0(c27_5_0, s28_5_0, s28_4_1, s28_6_0, c28_6_0);
	full_adder ad29_6_0(c28_5_0, s29_5_0, s29_4_1, s29_6_0, c29_6_0);
	full_adder ad30_6_0(c29_5_0, s30_5_0, s30_4_1, s30_6_0, c30_6_0);
	full_adder ad31_6_0(c30_5_0, s31_5_0, s31_5_1, s31_6_0, c31_6_0);
	full_adder ad32_6_0(c31_5_0, c31_5_1, s32_5_0, s32_6_0, c32_6_0);
	full_adder ad33_6_0(c32_5_0, c32_5_1, s33_5_0, s33_6_0, c33_6_0);
	full_adder ad34_6_0(c33_5_0, c33_5_1, s34_5_0, s34_6_0, c34_6_0);
	full_adder ad35_6_0(c34_5_0, c34_5_1, s35_5_0, s35_6_0, c35_6_0);
	full_adder ad36_6_0(c35_5_0, c35_5_1, s36_5_0, s36_6_0, c36_6_0);
	full_adder ad37_6_0(c36_5_0, c36_5_1, s37_5_0, s37_6_0, c37_6_0);
	full_adder ad38_6_0(c37_5_0, s38_5_0, s38_4_1, s38_6_0, c38_6_0);
	full_adder ad39_6_0(c38_5_0, s39_5_0, s39_4_1, s39_6_0, c39_6_0);
	full_adder ad40_6_0(c39_5_0, s40_5_0, s40_4_1, s40_6_0, c40_6_0);
	full_adder ad41_6_0(c40_5_0, s41_5_0, s41_4_1, s41_6_0, c41_6_0);
	full_adder ad42_6_0(c41_5_0, s42_5_0, s42_4_1, s42_6_0, c42_6_0);
	full_adder ad43_6_0(c42_5_0, s43_5_0, s43_4_1, s43_6_0, c43_6_0);
	full_adder ad44_6_0(c43_5_0, s44_5_0, s44_4_1, s44_6_0, c44_6_0);
	full_adder ad45_6_0(c44_5_0, s45_5_0, s45_3_1, s45_6_0, c45_6_0);
	half_adder ha46_6_0(c45_5_0, s46_5_0, s46_6_0, c46_6_0);
	half_adder ha47_6_0(c46_5_0, s47_5_0, s47_6_0, c47_6_0);
	half_adder ha48_6_0(c47_5_0, s48_5_0, s48_6_0, c48_6_0);
	half_adder ha49_6_0(c48_5_0, s49_5_0, s49_6_0, c49_6_0);
	half_adder ha50_6_0(c49_5_0, s50_5_0, s50_6_0, c50_6_0);
	half_adder ha51_6_0(c50_5_0, s51_5_0, s51_6_0, c51_6_0);
	half_adder ha52_6_0(c51_5_0, s52_5_0, s52_6_0, c52_6_0);
	half_adder ha53_6_0(c52_5_0, s53_5_0, s53_6_0, c53_6_0);
	half_adder ha54_6_0(c53_5_0, s54_5_0, s54_6_0, c54_6_0);
	half_adder ha55_6_0(c54_5_0, s55_5_0, s55_6_0, c55_6_0);
	half_adder ha56_6_0(c55_5_0, s56_5_0, s56_6_0, c56_6_0);
	half_adder ha57_6_0(c56_5_0, s57_5_0, s57_6_0, c57_6_0);
	half_adder ha58_6_0(c57_5_0, s58_5_0, s58_6_0, c58_6_0);
	half_adder ha59_6_0(c58_5_0, s59_5_0, s59_6_0, c59_6_0);
	half_adder ha60_6_0(c59_5_0, s60_5_0, s60_6_0, c60_6_0);
	half_adder ha61_6_0(c60_5_0, s61_5_0, s61_6_0, c61_6_0);
	half_adder ha62_6_0(c61_5_0, s62_5_0, s62_6_0, c62_6_0);
	half_adder ha63_6_0(c62_5_0, s63_5_0, s63_6_0, c63_6_0);

	half_adder ha8_7_0(c7_6_0, s8_6_0, s8_7_0, c8_7_0);
	half_adder ha9_7_0(c8_6_0, s9_6_0, s9_7_0, c9_7_0);
	half_adder ha10_7_0(c9_6_0, s10_6_0, s10_7_0, c10_7_0);
	half_adder ha11_7_0(c10_6_0, s11_6_0, s11_7_0, c11_7_0);
	half_adder ha12_7_0(c11_6_0, s12_6_0, s12_7_0, c12_7_0);
	half_adder ha13_7_0(c12_6_0, s13_6_0, s13_7_0, c13_7_0);
	half_adder ha14_7_0(c13_6_0, s14_6_0, s14_7_0, c14_7_0);
	half_adder ha15_7_0(c14_6_0, s15_6_0, s15_7_0, c15_7_0);
	half_adder ha16_7_0(c15_6_0, s16_6_0, s16_7_0, c16_7_0);
	half_adder ha17_7_0(c16_6_0, s17_6_0, s17_7_0, c17_7_0);
	half_adder ha18_7_0(c17_6_0, s18_6_0, s18_7_0, c18_7_0);
	half_adder ha19_7_0(c18_6_0, s19_6_0, s19_7_0, c19_7_0);
	half_adder ha20_7_0(c19_6_0, s20_6_0, s20_7_0, c20_7_0);
	half_adder ha21_7_0(c20_6_0, s21_6_0, s21_7_0, c21_7_0);
	half_adder ha22_7_0(c21_6_0, s22_6_0, s22_7_0, c22_7_0);
	half_adder ha23_7_0(c22_6_0, s23_6_0, s23_7_0, c23_7_0);
	half_adder ha24_7_0(c23_6_0, s24_6_0, s24_7_0, c24_7_0);
	half_adder ha25_7_0(c24_6_0, s25_6_0, s25_7_0, c25_7_0);
	half_adder ha26_7_0(c25_6_0, s26_6_0, s26_7_0, c26_7_0);
	half_adder ha27_7_0(c26_6_0, s27_6_0, s27_7_0, c27_7_0);
	half_adder ha28_7_0(c27_6_0, s28_6_0, s28_7_0, c28_7_0);
	half_adder ha29_7_0(c28_6_0, s29_6_0, s29_7_0, c29_7_0);
	half_adder ha30_7_0(c29_6_0, s30_6_0, s30_7_0, c30_7_0);
	half_adder ha31_7_0(c30_6_0, s31_6_0, s31_7_0, c31_7_0);
	full_adder ad32_7_0(c31_6_0, s32_6_0, s32_5_1, s32_7_0, c32_7_0);
	full_adder ad33_7_0(c32_6_0, s33_6_0, s33_5_1, s33_7_0, c33_7_0);
	full_adder ad34_7_0(c33_6_0, s34_6_0, s34_5_1, s34_7_0, c34_7_0);
	full_adder ad35_7_0(c34_6_0, s35_6_0, s35_5_1, s35_7_0, c35_7_0);
	full_adder ad36_7_0(c35_6_0, s36_6_0, s36_5_1, s36_7_0, c36_7_0);
	full_adder ad37_7_0(c36_6_0, s37_6_0, s37_4_1, s37_7_0, c37_7_0);
	half_adder ha38_7_0(c37_6_0, s38_6_0, s38_7_0, c38_7_0);
	half_adder ha39_7_0(c38_6_0, s39_6_0, s39_7_0, c39_7_0);
	half_adder ha40_7_0(c39_6_0, s40_6_0, s40_7_0, c40_7_0);
	half_adder ha41_7_0(c40_6_0, s41_6_0, s41_7_0, c41_7_0);
	half_adder ha42_7_0(c41_6_0, s42_6_0, s42_7_0, c42_7_0);
	half_adder ha43_7_0(c42_6_0, s43_6_0, s43_7_0, c43_7_0);
	half_adder ha44_7_0(c43_6_0, s44_6_0, s44_7_0, c44_7_0);
	half_adder ha45_7_0(c44_6_0, s45_6_0, s45_7_0, c45_7_0);
	half_adder ha46_7_0(c45_6_0, s46_6_0, s46_7_0, c46_7_0);
	half_adder ha47_7_0(c46_6_0, s47_6_0, s47_7_0, c47_7_0);
	half_adder ha48_7_0(c47_6_0, s48_6_0, s48_7_0, c48_7_0);
	half_adder ha49_7_0(c48_6_0, s49_6_0, s49_7_0, c49_7_0);
	half_adder ha50_7_0(c49_6_0, s50_6_0, s50_7_0, c50_7_0);
	half_adder ha51_7_0(c50_6_0, s51_6_0, s51_7_0, c51_7_0);
	half_adder ha52_7_0(c51_6_0, s52_6_0, s52_7_0, c52_7_0);
	half_adder ha53_7_0(c52_6_0, s53_6_0, s53_7_0, c53_7_0);
	half_adder ha54_7_0(c53_6_0, s54_6_0, s54_7_0, c54_7_0);
	half_adder ha55_7_0(c54_6_0, s55_6_0, s55_7_0, c55_7_0);
	half_adder ha56_7_0(c55_6_0, s56_6_0, s56_7_0, c56_7_0);
	half_adder ha57_7_0(c56_6_0, s57_6_0, s57_7_0, c57_7_0);
	half_adder ha58_7_0(c57_6_0, s58_6_0, s58_7_0, c58_7_0);
	half_adder ha59_7_0(c58_6_0, s59_6_0, s59_7_0, c59_7_0);
	half_adder ha60_7_0(c59_6_0, s60_6_0, s60_7_0, c60_7_0);
	half_adder ha61_7_0(c60_6_0, s61_6_0, s61_7_0, c61_7_0);
	half_adder ha62_7_0(c61_6_0, s62_6_0, s62_7_0, c62_7_0);
	half_adder ha63_7_0(c62_6_0, s63_6_0, s63_7_0, c63_7_0);


	assign x[0] = a0_0;
	assign x[1] = s1_0_0;
	assign x[2] = s2_1_0;
	assign x[3] = s3_2_0;
	assign x[4] = s4_3_0;
	assign x[5] = s5_4_0;
	assign x[6] = s6_5_0;
	assign x[7] = s7_6_0;
	assign x[8] = s8_7_0;
	assign x[9] = c8_7_0;
	assign x[10] = c9_7_0;
	assign x[11] = c10_7_0;
	assign x[12] = c11_7_0;
	assign x[13] = c12_7_0;
	assign x[14] = c13_7_0;
	assign x[15] = c14_7_0;
	assign x[16] = c15_7_0;
	assign x[17] = c16_7_0;
	assign x[18] = c17_7_0;
	assign x[19] = c18_7_0;
	assign x[20] = c19_7_0;
	assign x[21] = c20_7_0;
	assign x[22] = c21_7_0;
	assign x[23] = c22_7_0;
	assign x[24] = c23_7_0;
	assign x[25] = c24_7_0;
	assign x[26] = c25_7_0;
	assign x[27] = c26_7_0;
	assign x[28] = c27_7_0;
	assign x[29] = c28_7_0;
	assign x[30] = c29_7_0;
	assign x[31] = c30_7_0;
	assign x[32] = c31_7_0;
	assign x[33] = c32_7_0;
	assign x[34] = c33_7_0;
	assign x[35] = c34_7_0;
	assign x[36] = c35_7_0;
	assign x[37] = c36_7_0;
	assign x[38] = c37_7_0;
	assign x[39] = c38_7_0;
	assign x[40] = c39_7_0;
	assign x[41] = c40_7_0;
	assign x[42] = c41_7_0;
	assign x[43] = c42_7_0;
	assign x[44] = c43_7_0;
	assign x[45] = c44_7_0;
	assign x[46] = c45_7_0;
	assign x[47] = c46_7_0;
	assign x[48] = c47_7_0;
	assign x[49] = c48_7_0;
	assign x[50] = c49_7_0;
	assign x[51] = c50_7_0;
	assign x[52] = c51_7_0;
	assign x[53] = c52_7_0;
	assign x[54] = c53_7_0;
	assign x[55] = c54_7_0;
	assign x[56] = c55_7_0;
	assign x[57] = c56_7_0;
	assign x[58] = c57_7_0;
	assign x[59] = c58_7_0;
	assign x[60] = c59_7_0;
	assign x[61] = c60_7_0;
	assign x[62] = c61_7_0;
	assign x[63] = c62_7_0;
	assign y[0] = 1'b0;
	assign y[1] = 1'b0;
	assign y[2] = 1'b0;
	assign y[3] = 1'b0;
	assign y[4] = 1'b0;
	assign y[5] = 1'b0;
	assign y[6] = 1'b0;
	assign y[7] = 1'b0;
	assign y[8] = 1'b0;
	assign y[9] = s9_7_0;
	assign y[10] = s10_7_0;
	assign y[11] = s11_7_0;
	assign y[12] = s12_7_0;
	assign y[13] = s13_7_0;
	assign y[14] = s14_7_0;
	assign y[15] = s15_7_0;
	assign y[16] = s16_7_0;
	assign y[17] = s17_7_0;
	assign y[18] = s18_7_0;
	assign y[19] = s19_7_0;
	assign y[20] = s20_7_0;
	assign y[21] = s21_7_0;
	assign y[22] = s22_7_0;
	assign y[23] = s23_7_0;
	assign y[24] = s24_7_0;
	assign y[25] = s25_7_0;
	assign y[26] = s26_7_0;
	assign y[27] = s27_7_0;
	assign y[28] = s28_7_0;
	assign y[29] = s29_7_0;
	assign y[30] = s30_7_0;
	assign y[31] = s31_7_0;
	assign y[32] = s32_7_0;
	assign y[33] = s33_7_0;
	assign y[34] = s34_7_0;
	assign y[35] = s35_7_0;
	assign y[36] = s36_7_0;
	assign y[37] = s37_7_0;
	assign y[38] = s38_7_0;
	assign y[39] = s39_7_0;
	assign y[40] = s40_7_0;
	assign y[41] = s41_7_0;
	assign y[42] = s42_7_0;
	assign y[43] = s43_7_0;
	assign y[44] = s44_7_0;
	assign y[45] = s45_7_0;
	assign y[46] = s46_7_0;
	assign y[47] = s47_7_0;
	assign y[48] = s48_7_0;
	assign y[49] = s49_7_0;
	assign y[50] = s50_7_0;
	assign y[51] = s51_7_0;
	assign y[52] = s52_7_0;
	assign y[53] = s53_7_0;
	assign y[54] = s54_7_0;
	assign y[55] = s55_7_0;
	assign y[56] = s56_7_0;
	assign y[57] = s57_7_0;
	assign y[58] = s58_7_0;
	assign y[59] = s59_7_0;
	assign y[60] = s60_7_0;
	assign y[61] = s61_7_0;
	assign y[62] = s62_7_0;
	assign y[63] = s63_7_0;

	carry_select_32 cs32_0(1'b0, x[31:0], y[31:0], cout, product);
	
	carry_select_32 cs32_1a(1'b0, x[63:32], y[63:32], cout_a, upperbits_a);
	carry_select_32 cs32_1b(1'b1, x[63:32], y[63:32], cout_b, upperbits_b);
	
	mux_2 cs_mux(cout, upperbits_a, upperbits_b, upperbits);
	
	xor xo0(xo_0, upperbits[0], upperbits[16]);
	xor xo1(xo_1, upperbits[1], upperbits[17]);
	xor xo2(xo_2, upperbits[2], upperbits[18]);
	xor xo3(xo_3, upperbits[3], upperbits[19]);
	xor xo4(xo_4, upperbits[4], upperbits[20]);
	xor xo5(xo_5, upperbits[5], upperbits[21]);
	xor xo6(xo_6, upperbits[6], upperbits[22]);
	xor xo7(xo_7, upperbits[7], upperbits[23]);
	xor xo8(xo_8, upperbits[8], upperbits[24]);
	xor xo9(xo_9, upperbits[9], upperbits[25]);
	xor xo10(xo_10, upperbits[10], upperbits[26]);
	xor xo11(xo_11, upperbits[11], upperbits[27]);
	xor xo12(xo_12, upperbits[12], upperbits[28]);
	xor xo13(xo_13, upperbits[13], upperbits[29]);
	xor xo14(xo_14, upperbits[14], upperbits[30]);
	xor xo15(xo_15, upperbits[15], upperbits[31]);
	
	or o0(o_0, xo_0, xo_1, xo_2, xo_3);
	or o1(o_1, xo_4, xo_5, xo_6, xo_7);
	or o2(o_2, xo_8, xo_9, xo_10, xo_11);
	or o3(o_3, xo_12, xo_13, xo_14, xo_15);
	
	or o4(o_4, o_0, o_1, o_2, o_3); //checks to see if all upper bits are the same; should be 0
	
	not n0(n_0, o_4); //should be 1 if all upper bits are same
	
	xnor xno0(xno_0, upperbits[0], product[31]); //check to see if upper bits and sign extension are the same, 1 if they are
	
	and a0(n_overflow, n_0, xno_0); //if all upper bits are the same AND they're the same as the top bit we're good
	
	not n1(overflow, n_overflow);

endmodule
