module mips_tb()


endmodule 